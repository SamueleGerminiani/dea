
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_myproject.layer2_out_V_U.if_read & AESL_inst_myproject.layer2_out_V_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_myproject.layer2_out_V_U.if_write & AESL_inst_myproject.layer2_out_V_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = 0;
    assign fifo_intf_1.fifo_wr_block = 0;
    assign fifo_intf_1.finish = finish;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_myproject.layer2_out_V_1_U.if_read & AESL_inst_myproject.layer2_out_V_1_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_myproject.layer2_out_V_1_U.if_write & AESL_inst_myproject.layer2_out_V_1_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = 0;
    assign fifo_intf_2.fifo_wr_block = 0;
    assign fifo_intf_2.finish = finish;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_myproject.layer2_out_V_2_U.if_read & AESL_inst_myproject.layer2_out_V_2_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_myproject.layer2_out_V_2_U.if_write & AESL_inst_myproject.layer2_out_V_2_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = 0;
    assign fifo_intf_3.fifo_wr_block = 0;
    assign fifo_intf_3.finish = finish;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_myproject.layer2_out_V_3_U.if_read & AESL_inst_myproject.layer2_out_V_3_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_myproject.layer2_out_V_3_U.if_write & AESL_inst_myproject.layer2_out_V_3_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = 0;
    assign fifo_intf_4.fifo_wr_block = 0;
    assign fifo_intf_4.finish = finish;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_myproject.layer2_out_V_4_U.if_read & AESL_inst_myproject.layer2_out_V_4_U.if_empty_n;
    assign fifo_intf_5.wr_en = AESL_inst_myproject.layer2_out_V_4_U.if_write & AESL_inst_myproject.layer2_out_V_4_U.if_full_n;
    assign fifo_intf_5.fifo_rd_block = 0;
    assign fifo_intf_5.fifo_wr_block = 0;
    assign fifo_intf_5.finish = finish;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_myproject.layer2_out_V_5_U.if_read & AESL_inst_myproject.layer2_out_V_5_U.if_empty_n;
    assign fifo_intf_6.wr_en = AESL_inst_myproject.layer2_out_V_5_U.if_write & AESL_inst_myproject.layer2_out_V_5_U.if_full_n;
    assign fifo_intf_6.fifo_rd_block = 0;
    assign fifo_intf_6.fifo_wr_block = 0;
    assign fifo_intf_6.finish = finish;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_myproject.layer2_out_V_6_U.if_read & AESL_inst_myproject.layer2_out_V_6_U.if_empty_n;
    assign fifo_intf_7.wr_en = AESL_inst_myproject.layer2_out_V_6_U.if_write & AESL_inst_myproject.layer2_out_V_6_U.if_full_n;
    assign fifo_intf_7.fifo_rd_block = 0;
    assign fifo_intf_7.fifo_wr_block = 0;
    assign fifo_intf_7.finish = finish;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_myproject.layer2_out_V_7_U.if_read & AESL_inst_myproject.layer2_out_V_7_U.if_empty_n;
    assign fifo_intf_8.wr_en = AESL_inst_myproject.layer2_out_V_7_U.if_write & AESL_inst_myproject.layer2_out_V_7_U.if_full_n;
    assign fifo_intf_8.fifo_rd_block = 0;
    assign fifo_intf_8.fifo_wr_block = 0;
    assign fifo_intf_8.finish = finish;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_myproject.layer2_out_V_8_U.if_read & AESL_inst_myproject.layer2_out_V_8_U.if_empty_n;
    assign fifo_intf_9.wr_en = AESL_inst_myproject.layer2_out_V_8_U.if_write & AESL_inst_myproject.layer2_out_V_8_U.if_full_n;
    assign fifo_intf_9.fifo_rd_block = 0;
    assign fifo_intf_9.fifo_wr_block = 0;
    assign fifo_intf_9.finish = finish;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_myproject.layer2_out_V_9_U.if_read & AESL_inst_myproject.layer2_out_V_9_U.if_empty_n;
    assign fifo_intf_10.wr_en = AESL_inst_myproject.layer2_out_V_9_U.if_write & AESL_inst_myproject.layer2_out_V_9_U.if_full_n;
    assign fifo_intf_10.fifo_rd_block = 0;
    assign fifo_intf_10.fifo_wr_block = 0;
    assign fifo_intf_10.finish = finish;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_myproject.layer2_out_V_10_U.if_read & AESL_inst_myproject.layer2_out_V_10_U.if_empty_n;
    assign fifo_intf_11.wr_en = AESL_inst_myproject.layer2_out_V_10_U.if_write & AESL_inst_myproject.layer2_out_V_10_U.if_full_n;
    assign fifo_intf_11.fifo_rd_block = 0;
    assign fifo_intf_11.fifo_wr_block = 0;
    assign fifo_intf_11.finish = finish;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_myproject.layer2_out_V_11_U.if_read & AESL_inst_myproject.layer2_out_V_11_U.if_empty_n;
    assign fifo_intf_12.wr_en = AESL_inst_myproject.layer2_out_V_11_U.if_write & AESL_inst_myproject.layer2_out_V_11_U.if_full_n;
    assign fifo_intf_12.fifo_rd_block = 0;
    assign fifo_intf_12.fifo_wr_block = 0;
    assign fifo_intf_12.finish = finish;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_myproject.layer2_out_V_12_U.if_read & AESL_inst_myproject.layer2_out_V_12_U.if_empty_n;
    assign fifo_intf_13.wr_en = AESL_inst_myproject.layer2_out_V_12_U.if_write & AESL_inst_myproject.layer2_out_V_12_U.if_full_n;
    assign fifo_intf_13.fifo_rd_block = 0;
    assign fifo_intf_13.fifo_wr_block = 0;
    assign fifo_intf_13.finish = finish;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_myproject.layer2_out_V_13_U.if_read & AESL_inst_myproject.layer2_out_V_13_U.if_empty_n;
    assign fifo_intf_14.wr_en = AESL_inst_myproject.layer2_out_V_13_U.if_write & AESL_inst_myproject.layer2_out_V_13_U.if_full_n;
    assign fifo_intf_14.fifo_rd_block = 0;
    assign fifo_intf_14.fifo_wr_block = 0;
    assign fifo_intf_14.finish = finish;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_myproject.layer2_out_V_14_U.if_read & AESL_inst_myproject.layer2_out_V_14_U.if_empty_n;
    assign fifo_intf_15.wr_en = AESL_inst_myproject.layer2_out_V_14_U.if_write & AESL_inst_myproject.layer2_out_V_14_U.if_full_n;
    assign fifo_intf_15.fifo_rd_block = 0;
    assign fifo_intf_15.fifo_wr_block = 0;
    assign fifo_intf_15.finish = finish;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_myproject.layer2_out_V_15_U.if_read & AESL_inst_myproject.layer2_out_V_15_U.if_empty_n;
    assign fifo_intf_16.wr_en = AESL_inst_myproject.layer2_out_V_15_U.if_write & AESL_inst_myproject.layer2_out_V_15_U.if_full_n;
    assign fifo_intf_16.fifo_rd_block = 0;
    assign fifo_intf_16.fifo_wr_block = 0;
    assign fifo_intf_16.finish = finish;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_myproject.layer2_out_V_16_U.if_read & AESL_inst_myproject.layer2_out_V_16_U.if_empty_n;
    assign fifo_intf_17.wr_en = AESL_inst_myproject.layer2_out_V_16_U.if_write & AESL_inst_myproject.layer2_out_V_16_U.if_full_n;
    assign fifo_intf_17.fifo_rd_block = 0;
    assign fifo_intf_17.fifo_wr_block = 0;
    assign fifo_intf_17.finish = finish;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;
    df_fifo_intf fifo_intf_18(clock,reset);
    assign fifo_intf_18.rd_en = AESL_inst_myproject.layer2_out_V_17_U.if_read & AESL_inst_myproject.layer2_out_V_17_U.if_empty_n;
    assign fifo_intf_18.wr_en = AESL_inst_myproject.layer2_out_V_17_U.if_write & AESL_inst_myproject.layer2_out_V_17_U.if_full_n;
    assign fifo_intf_18.fifo_rd_block = 0;
    assign fifo_intf_18.fifo_wr_block = 0;
    assign fifo_intf_18.finish = finish;
    csv_file_dump fifo_csv_dumper_18;
    csv_file_dump cstatus_csv_dumper_18;
    df_fifo_monitor fifo_monitor_18;
    df_fifo_intf fifo_intf_19(clock,reset);
    assign fifo_intf_19.rd_en = AESL_inst_myproject.layer2_out_V_18_U.if_read & AESL_inst_myproject.layer2_out_V_18_U.if_empty_n;
    assign fifo_intf_19.wr_en = AESL_inst_myproject.layer2_out_V_18_U.if_write & AESL_inst_myproject.layer2_out_V_18_U.if_full_n;
    assign fifo_intf_19.fifo_rd_block = 0;
    assign fifo_intf_19.fifo_wr_block = 0;
    assign fifo_intf_19.finish = finish;
    csv_file_dump fifo_csv_dumper_19;
    csv_file_dump cstatus_csv_dumper_19;
    df_fifo_monitor fifo_monitor_19;
    df_fifo_intf fifo_intf_20(clock,reset);
    assign fifo_intf_20.rd_en = AESL_inst_myproject.layer2_out_V_19_U.if_read & AESL_inst_myproject.layer2_out_V_19_U.if_empty_n;
    assign fifo_intf_20.wr_en = AESL_inst_myproject.layer2_out_V_19_U.if_write & AESL_inst_myproject.layer2_out_V_19_U.if_full_n;
    assign fifo_intf_20.fifo_rd_block = 0;
    assign fifo_intf_20.fifo_wr_block = 0;
    assign fifo_intf_20.finish = finish;
    csv_file_dump fifo_csv_dumper_20;
    csv_file_dump cstatus_csv_dumper_20;
    df_fifo_monitor fifo_monitor_20;
    df_fifo_intf fifo_intf_21(clock,reset);
    assign fifo_intf_21.rd_en = AESL_inst_myproject.layer2_out_V_20_U.if_read & AESL_inst_myproject.layer2_out_V_20_U.if_empty_n;
    assign fifo_intf_21.wr_en = AESL_inst_myproject.layer2_out_V_20_U.if_write & AESL_inst_myproject.layer2_out_V_20_U.if_full_n;
    assign fifo_intf_21.fifo_rd_block = 0;
    assign fifo_intf_21.fifo_wr_block = 0;
    assign fifo_intf_21.finish = finish;
    csv_file_dump fifo_csv_dumper_21;
    csv_file_dump cstatus_csv_dumper_21;
    df_fifo_monitor fifo_monitor_21;
    df_fifo_intf fifo_intf_22(clock,reset);
    assign fifo_intf_22.rd_en = AESL_inst_myproject.layer2_out_V_21_U.if_read & AESL_inst_myproject.layer2_out_V_21_U.if_empty_n;
    assign fifo_intf_22.wr_en = AESL_inst_myproject.layer2_out_V_21_U.if_write & AESL_inst_myproject.layer2_out_V_21_U.if_full_n;
    assign fifo_intf_22.fifo_rd_block = 0;
    assign fifo_intf_22.fifo_wr_block = 0;
    assign fifo_intf_22.finish = finish;
    csv_file_dump fifo_csv_dumper_22;
    csv_file_dump cstatus_csv_dumper_22;
    df_fifo_monitor fifo_monitor_22;
    df_fifo_intf fifo_intf_23(clock,reset);
    assign fifo_intf_23.rd_en = AESL_inst_myproject.layer2_out_V_22_U.if_read & AESL_inst_myproject.layer2_out_V_22_U.if_empty_n;
    assign fifo_intf_23.wr_en = AESL_inst_myproject.layer2_out_V_22_U.if_write & AESL_inst_myproject.layer2_out_V_22_U.if_full_n;
    assign fifo_intf_23.fifo_rd_block = 0;
    assign fifo_intf_23.fifo_wr_block = 0;
    assign fifo_intf_23.finish = finish;
    csv_file_dump fifo_csv_dumper_23;
    csv_file_dump cstatus_csv_dumper_23;
    df_fifo_monitor fifo_monitor_23;
    df_fifo_intf fifo_intf_24(clock,reset);
    assign fifo_intf_24.rd_en = AESL_inst_myproject.layer2_out_V_23_U.if_read & AESL_inst_myproject.layer2_out_V_23_U.if_empty_n;
    assign fifo_intf_24.wr_en = AESL_inst_myproject.layer2_out_V_23_U.if_write & AESL_inst_myproject.layer2_out_V_23_U.if_full_n;
    assign fifo_intf_24.fifo_rd_block = 0;
    assign fifo_intf_24.fifo_wr_block = 0;
    assign fifo_intf_24.finish = finish;
    csv_file_dump fifo_csv_dumper_24;
    csv_file_dump cstatus_csv_dumper_24;
    df_fifo_monitor fifo_monitor_24;
    df_fifo_intf fifo_intf_25(clock,reset);
    assign fifo_intf_25.rd_en = AESL_inst_myproject.layer2_out_V_24_U.if_read & AESL_inst_myproject.layer2_out_V_24_U.if_empty_n;
    assign fifo_intf_25.wr_en = AESL_inst_myproject.layer2_out_V_24_U.if_write & AESL_inst_myproject.layer2_out_V_24_U.if_full_n;
    assign fifo_intf_25.fifo_rd_block = 0;
    assign fifo_intf_25.fifo_wr_block = 0;
    assign fifo_intf_25.finish = finish;
    csv_file_dump fifo_csv_dumper_25;
    csv_file_dump cstatus_csv_dumper_25;
    df_fifo_monitor fifo_monitor_25;
    df_fifo_intf fifo_intf_26(clock,reset);
    assign fifo_intf_26.rd_en = AESL_inst_myproject.layer2_out_V_25_U.if_read & AESL_inst_myproject.layer2_out_V_25_U.if_empty_n;
    assign fifo_intf_26.wr_en = AESL_inst_myproject.layer2_out_V_25_U.if_write & AESL_inst_myproject.layer2_out_V_25_U.if_full_n;
    assign fifo_intf_26.fifo_rd_block = 0;
    assign fifo_intf_26.fifo_wr_block = 0;
    assign fifo_intf_26.finish = finish;
    csv_file_dump fifo_csv_dumper_26;
    csv_file_dump cstatus_csv_dumper_26;
    df_fifo_monitor fifo_monitor_26;
    df_fifo_intf fifo_intf_27(clock,reset);
    assign fifo_intf_27.rd_en = AESL_inst_myproject.layer2_out_V_26_U.if_read & AESL_inst_myproject.layer2_out_V_26_U.if_empty_n;
    assign fifo_intf_27.wr_en = AESL_inst_myproject.layer2_out_V_26_U.if_write & AESL_inst_myproject.layer2_out_V_26_U.if_full_n;
    assign fifo_intf_27.fifo_rd_block = 0;
    assign fifo_intf_27.fifo_wr_block = 0;
    assign fifo_intf_27.finish = finish;
    csv_file_dump fifo_csv_dumper_27;
    csv_file_dump cstatus_csv_dumper_27;
    df_fifo_monitor fifo_monitor_27;
    df_fifo_intf fifo_intf_28(clock,reset);
    assign fifo_intf_28.rd_en = AESL_inst_myproject.layer2_out_V_27_U.if_read & AESL_inst_myproject.layer2_out_V_27_U.if_empty_n;
    assign fifo_intf_28.wr_en = AESL_inst_myproject.layer2_out_V_27_U.if_write & AESL_inst_myproject.layer2_out_V_27_U.if_full_n;
    assign fifo_intf_28.fifo_rd_block = 0;
    assign fifo_intf_28.fifo_wr_block = 0;
    assign fifo_intf_28.finish = finish;
    csv_file_dump fifo_csv_dumper_28;
    csv_file_dump cstatus_csv_dumper_28;
    df_fifo_monitor fifo_monitor_28;
    df_fifo_intf fifo_intf_29(clock,reset);
    assign fifo_intf_29.rd_en = AESL_inst_myproject.layer2_out_V_28_U.if_read & AESL_inst_myproject.layer2_out_V_28_U.if_empty_n;
    assign fifo_intf_29.wr_en = AESL_inst_myproject.layer2_out_V_28_U.if_write & AESL_inst_myproject.layer2_out_V_28_U.if_full_n;
    assign fifo_intf_29.fifo_rd_block = 0;
    assign fifo_intf_29.fifo_wr_block = 0;
    assign fifo_intf_29.finish = finish;
    csv_file_dump fifo_csv_dumper_29;
    csv_file_dump cstatus_csv_dumper_29;
    df_fifo_monitor fifo_monitor_29;
    df_fifo_intf fifo_intf_30(clock,reset);
    assign fifo_intf_30.rd_en = AESL_inst_myproject.layer2_out_V_29_U.if_read & AESL_inst_myproject.layer2_out_V_29_U.if_empty_n;
    assign fifo_intf_30.wr_en = AESL_inst_myproject.layer2_out_V_29_U.if_write & AESL_inst_myproject.layer2_out_V_29_U.if_full_n;
    assign fifo_intf_30.fifo_rd_block = 0;
    assign fifo_intf_30.fifo_wr_block = 0;
    assign fifo_intf_30.finish = finish;
    csv_file_dump fifo_csv_dumper_30;
    csv_file_dump cstatus_csv_dumper_30;
    df_fifo_monitor fifo_monitor_30;
    df_fifo_intf fifo_intf_31(clock,reset);
    assign fifo_intf_31.rd_en = AESL_inst_myproject.layer2_out_V_30_U.if_read & AESL_inst_myproject.layer2_out_V_30_U.if_empty_n;
    assign fifo_intf_31.wr_en = AESL_inst_myproject.layer2_out_V_30_U.if_write & AESL_inst_myproject.layer2_out_V_30_U.if_full_n;
    assign fifo_intf_31.fifo_rd_block = 0;
    assign fifo_intf_31.fifo_wr_block = 0;
    assign fifo_intf_31.finish = finish;
    csv_file_dump fifo_csv_dumper_31;
    csv_file_dump cstatus_csv_dumper_31;
    df_fifo_monitor fifo_monitor_31;
    df_fifo_intf fifo_intf_32(clock,reset);
    assign fifo_intf_32.rd_en = AESL_inst_myproject.layer2_out_V_31_U.if_read & AESL_inst_myproject.layer2_out_V_31_U.if_empty_n;
    assign fifo_intf_32.wr_en = AESL_inst_myproject.layer2_out_V_31_U.if_write & AESL_inst_myproject.layer2_out_V_31_U.if_full_n;
    assign fifo_intf_32.fifo_rd_block = 0;
    assign fifo_intf_32.fifo_wr_block = 0;
    assign fifo_intf_32.finish = finish;
    csv_file_dump fifo_csv_dumper_32;
    csv_file_dump cstatus_csv_dumper_32;
    df_fifo_monitor fifo_monitor_32;
    df_fifo_intf fifo_intf_33(clock,reset);
    assign fifo_intf_33.rd_en = AESL_inst_myproject.layer2_out_V_32_U.if_read & AESL_inst_myproject.layer2_out_V_32_U.if_empty_n;
    assign fifo_intf_33.wr_en = AESL_inst_myproject.layer2_out_V_32_U.if_write & AESL_inst_myproject.layer2_out_V_32_U.if_full_n;
    assign fifo_intf_33.fifo_rd_block = 0;
    assign fifo_intf_33.fifo_wr_block = 0;
    assign fifo_intf_33.finish = finish;
    csv_file_dump fifo_csv_dumper_33;
    csv_file_dump cstatus_csv_dumper_33;
    df_fifo_monitor fifo_monitor_33;
    df_fifo_intf fifo_intf_34(clock,reset);
    assign fifo_intf_34.rd_en = AESL_inst_myproject.layer2_out_V_33_U.if_read & AESL_inst_myproject.layer2_out_V_33_U.if_empty_n;
    assign fifo_intf_34.wr_en = AESL_inst_myproject.layer2_out_V_33_U.if_write & AESL_inst_myproject.layer2_out_V_33_U.if_full_n;
    assign fifo_intf_34.fifo_rd_block = 0;
    assign fifo_intf_34.fifo_wr_block = 0;
    assign fifo_intf_34.finish = finish;
    csv_file_dump fifo_csv_dumper_34;
    csv_file_dump cstatus_csv_dumper_34;
    df_fifo_monitor fifo_monitor_34;
    df_fifo_intf fifo_intf_35(clock,reset);
    assign fifo_intf_35.rd_en = AESL_inst_myproject.layer2_out_V_34_U.if_read & AESL_inst_myproject.layer2_out_V_34_U.if_empty_n;
    assign fifo_intf_35.wr_en = AESL_inst_myproject.layer2_out_V_34_U.if_write & AESL_inst_myproject.layer2_out_V_34_U.if_full_n;
    assign fifo_intf_35.fifo_rd_block = 0;
    assign fifo_intf_35.fifo_wr_block = 0;
    assign fifo_intf_35.finish = finish;
    csv_file_dump fifo_csv_dumper_35;
    csv_file_dump cstatus_csv_dumper_35;
    df_fifo_monitor fifo_monitor_35;
    df_fifo_intf fifo_intf_36(clock,reset);
    assign fifo_intf_36.rd_en = AESL_inst_myproject.layer2_out_V_35_U.if_read & AESL_inst_myproject.layer2_out_V_35_U.if_empty_n;
    assign fifo_intf_36.wr_en = AESL_inst_myproject.layer2_out_V_35_U.if_write & AESL_inst_myproject.layer2_out_V_35_U.if_full_n;
    assign fifo_intf_36.fifo_rd_block = 0;
    assign fifo_intf_36.fifo_wr_block = 0;
    assign fifo_intf_36.finish = finish;
    csv_file_dump fifo_csv_dumper_36;
    csv_file_dump cstatus_csv_dumper_36;
    df_fifo_monitor fifo_monitor_36;
    df_fifo_intf fifo_intf_37(clock,reset);
    assign fifo_intf_37.rd_en = AESL_inst_myproject.layer2_out_V_36_U.if_read & AESL_inst_myproject.layer2_out_V_36_U.if_empty_n;
    assign fifo_intf_37.wr_en = AESL_inst_myproject.layer2_out_V_36_U.if_write & AESL_inst_myproject.layer2_out_V_36_U.if_full_n;
    assign fifo_intf_37.fifo_rd_block = 0;
    assign fifo_intf_37.fifo_wr_block = 0;
    assign fifo_intf_37.finish = finish;
    csv_file_dump fifo_csv_dumper_37;
    csv_file_dump cstatus_csv_dumper_37;
    df_fifo_monitor fifo_monitor_37;
    df_fifo_intf fifo_intf_38(clock,reset);
    assign fifo_intf_38.rd_en = AESL_inst_myproject.layer2_out_V_37_U.if_read & AESL_inst_myproject.layer2_out_V_37_U.if_empty_n;
    assign fifo_intf_38.wr_en = AESL_inst_myproject.layer2_out_V_37_U.if_write & AESL_inst_myproject.layer2_out_V_37_U.if_full_n;
    assign fifo_intf_38.fifo_rd_block = 0;
    assign fifo_intf_38.fifo_wr_block = 0;
    assign fifo_intf_38.finish = finish;
    csv_file_dump fifo_csv_dumper_38;
    csv_file_dump cstatus_csv_dumper_38;
    df_fifo_monitor fifo_monitor_38;
    df_fifo_intf fifo_intf_39(clock,reset);
    assign fifo_intf_39.rd_en = AESL_inst_myproject.layer2_out_V_38_U.if_read & AESL_inst_myproject.layer2_out_V_38_U.if_empty_n;
    assign fifo_intf_39.wr_en = AESL_inst_myproject.layer2_out_V_38_U.if_write & AESL_inst_myproject.layer2_out_V_38_U.if_full_n;
    assign fifo_intf_39.fifo_rd_block = 0;
    assign fifo_intf_39.fifo_wr_block = 0;
    assign fifo_intf_39.finish = finish;
    csv_file_dump fifo_csv_dumper_39;
    csv_file_dump cstatus_csv_dumper_39;
    df_fifo_monitor fifo_monitor_39;
    df_fifo_intf fifo_intf_40(clock,reset);
    assign fifo_intf_40.rd_en = AESL_inst_myproject.layer2_out_V_39_U.if_read & AESL_inst_myproject.layer2_out_V_39_U.if_empty_n;
    assign fifo_intf_40.wr_en = AESL_inst_myproject.layer2_out_V_39_U.if_write & AESL_inst_myproject.layer2_out_V_39_U.if_full_n;
    assign fifo_intf_40.fifo_rd_block = 0;
    assign fifo_intf_40.fifo_wr_block = 0;
    assign fifo_intf_40.finish = finish;
    csv_file_dump fifo_csv_dumper_40;
    csv_file_dump cstatus_csv_dumper_40;
    df_fifo_monitor fifo_monitor_40;
    df_fifo_intf fifo_intf_41(clock,reset);
    assign fifo_intf_41.rd_en = AESL_inst_myproject.layer2_out_V_40_U.if_read & AESL_inst_myproject.layer2_out_V_40_U.if_empty_n;
    assign fifo_intf_41.wr_en = AESL_inst_myproject.layer2_out_V_40_U.if_write & AESL_inst_myproject.layer2_out_V_40_U.if_full_n;
    assign fifo_intf_41.fifo_rd_block = 0;
    assign fifo_intf_41.fifo_wr_block = 0;
    assign fifo_intf_41.finish = finish;
    csv_file_dump fifo_csv_dumper_41;
    csv_file_dump cstatus_csv_dumper_41;
    df_fifo_monitor fifo_monitor_41;
    df_fifo_intf fifo_intf_42(clock,reset);
    assign fifo_intf_42.rd_en = AESL_inst_myproject.layer2_out_V_41_U.if_read & AESL_inst_myproject.layer2_out_V_41_U.if_empty_n;
    assign fifo_intf_42.wr_en = AESL_inst_myproject.layer2_out_V_41_U.if_write & AESL_inst_myproject.layer2_out_V_41_U.if_full_n;
    assign fifo_intf_42.fifo_rd_block = 0;
    assign fifo_intf_42.fifo_wr_block = 0;
    assign fifo_intf_42.finish = finish;
    csv_file_dump fifo_csv_dumper_42;
    csv_file_dump cstatus_csv_dumper_42;
    df_fifo_monitor fifo_monitor_42;
    df_fifo_intf fifo_intf_43(clock,reset);
    assign fifo_intf_43.rd_en = AESL_inst_myproject.layer2_out_V_42_U.if_read & AESL_inst_myproject.layer2_out_V_42_U.if_empty_n;
    assign fifo_intf_43.wr_en = AESL_inst_myproject.layer2_out_V_42_U.if_write & AESL_inst_myproject.layer2_out_V_42_U.if_full_n;
    assign fifo_intf_43.fifo_rd_block = 0;
    assign fifo_intf_43.fifo_wr_block = 0;
    assign fifo_intf_43.finish = finish;
    csv_file_dump fifo_csv_dumper_43;
    csv_file_dump cstatus_csv_dumper_43;
    df_fifo_monitor fifo_monitor_43;
    df_fifo_intf fifo_intf_44(clock,reset);
    assign fifo_intf_44.rd_en = AESL_inst_myproject.layer2_out_V_43_U.if_read & AESL_inst_myproject.layer2_out_V_43_U.if_empty_n;
    assign fifo_intf_44.wr_en = AESL_inst_myproject.layer2_out_V_43_U.if_write & AESL_inst_myproject.layer2_out_V_43_U.if_full_n;
    assign fifo_intf_44.fifo_rd_block = 0;
    assign fifo_intf_44.fifo_wr_block = 0;
    assign fifo_intf_44.finish = finish;
    csv_file_dump fifo_csv_dumper_44;
    csv_file_dump cstatus_csv_dumper_44;
    df_fifo_monitor fifo_monitor_44;
    df_fifo_intf fifo_intf_45(clock,reset);
    assign fifo_intf_45.rd_en = AESL_inst_myproject.layer2_out_V_44_U.if_read & AESL_inst_myproject.layer2_out_V_44_U.if_empty_n;
    assign fifo_intf_45.wr_en = AESL_inst_myproject.layer2_out_V_44_U.if_write & AESL_inst_myproject.layer2_out_V_44_U.if_full_n;
    assign fifo_intf_45.fifo_rd_block = 0;
    assign fifo_intf_45.fifo_wr_block = 0;
    assign fifo_intf_45.finish = finish;
    csv_file_dump fifo_csv_dumper_45;
    csv_file_dump cstatus_csv_dumper_45;
    df_fifo_monitor fifo_monitor_45;
    df_fifo_intf fifo_intf_46(clock,reset);
    assign fifo_intf_46.rd_en = AESL_inst_myproject.layer2_out_V_45_U.if_read & AESL_inst_myproject.layer2_out_V_45_U.if_empty_n;
    assign fifo_intf_46.wr_en = AESL_inst_myproject.layer2_out_V_45_U.if_write & AESL_inst_myproject.layer2_out_V_45_U.if_full_n;
    assign fifo_intf_46.fifo_rd_block = 0;
    assign fifo_intf_46.fifo_wr_block = 0;
    assign fifo_intf_46.finish = finish;
    csv_file_dump fifo_csv_dumper_46;
    csv_file_dump cstatus_csv_dumper_46;
    df_fifo_monitor fifo_monitor_46;
    df_fifo_intf fifo_intf_47(clock,reset);
    assign fifo_intf_47.rd_en = AESL_inst_myproject.layer2_out_V_46_U.if_read & AESL_inst_myproject.layer2_out_V_46_U.if_empty_n;
    assign fifo_intf_47.wr_en = AESL_inst_myproject.layer2_out_V_46_U.if_write & AESL_inst_myproject.layer2_out_V_46_U.if_full_n;
    assign fifo_intf_47.fifo_rd_block = 0;
    assign fifo_intf_47.fifo_wr_block = 0;
    assign fifo_intf_47.finish = finish;
    csv_file_dump fifo_csv_dumper_47;
    csv_file_dump cstatus_csv_dumper_47;
    df_fifo_monitor fifo_monitor_47;
    df_fifo_intf fifo_intf_48(clock,reset);
    assign fifo_intf_48.rd_en = AESL_inst_myproject.layer2_out_V_47_U.if_read & AESL_inst_myproject.layer2_out_V_47_U.if_empty_n;
    assign fifo_intf_48.wr_en = AESL_inst_myproject.layer2_out_V_47_U.if_write & AESL_inst_myproject.layer2_out_V_47_U.if_full_n;
    assign fifo_intf_48.fifo_rd_block = 0;
    assign fifo_intf_48.fifo_wr_block = 0;
    assign fifo_intf_48.finish = finish;
    csv_file_dump fifo_csv_dumper_48;
    csv_file_dump cstatus_csv_dumper_48;
    df_fifo_monitor fifo_monitor_48;
    df_fifo_intf fifo_intf_49(clock,reset);
    assign fifo_intf_49.rd_en = AESL_inst_myproject.layer2_out_V_48_U.if_read & AESL_inst_myproject.layer2_out_V_48_U.if_empty_n;
    assign fifo_intf_49.wr_en = AESL_inst_myproject.layer2_out_V_48_U.if_write & AESL_inst_myproject.layer2_out_V_48_U.if_full_n;
    assign fifo_intf_49.fifo_rd_block = 0;
    assign fifo_intf_49.fifo_wr_block = 0;
    assign fifo_intf_49.finish = finish;
    csv_file_dump fifo_csv_dumper_49;
    csv_file_dump cstatus_csv_dumper_49;
    df_fifo_monitor fifo_monitor_49;
    df_fifo_intf fifo_intf_50(clock,reset);
    assign fifo_intf_50.rd_en = AESL_inst_myproject.layer2_out_V_49_U.if_read & AESL_inst_myproject.layer2_out_V_49_U.if_empty_n;
    assign fifo_intf_50.wr_en = AESL_inst_myproject.layer2_out_V_49_U.if_write & AESL_inst_myproject.layer2_out_V_49_U.if_full_n;
    assign fifo_intf_50.fifo_rd_block = 0;
    assign fifo_intf_50.fifo_wr_block = 0;
    assign fifo_intf_50.finish = finish;
    csv_file_dump fifo_csv_dumper_50;
    csv_file_dump cstatus_csv_dumper_50;
    df_fifo_monitor fifo_monitor_50;
    df_fifo_intf fifo_intf_51(clock,reset);
    assign fifo_intf_51.rd_en = AESL_inst_myproject.layer4_out_V_U.if_read & AESL_inst_myproject.layer4_out_V_U.if_empty_n;
    assign fifo_intf_51.wr_en = AESL_inst_myproject.layer4_out_V_U.if_write & AESL_inst_myproject.layer4_out_V_U.if_full_n;
    assign fifo_intf_51.fifo_rd_block = 0;
    assign fifo_intf_51.fifo_wr_block = 0;
    assign fifo_intf_51.finish = finish;
    csv_file_dump fifo_csv_dumper_51;
    csv_file_dump cstatus_csv_dumper_51;
    df_fifo_monitor fifo_monitor_51;
    df_fifo_intf fifo_intf_52(clock,reset);
    assign fifo_intf_52.rd_en = AESL_inst_myproject.layer4_out_V_1_U.if_read & AESL_inst_myproject.layer4_out_V_1_U.if_empty_n;
    assign fifo_intf_52.wr_en = AESL_inst_myproject.layer4_out_V_1_U.if_write & AESL_inst_myproject.layer4_out_V_1_U.if_full_n;
    assign fifo_intf_52.fifo_rd_block = 0;
    assign fifo_intf_52.fifo_wr_block = 0;
    assign fifo_intf_52.finish = finish;
    csv_file_dump fifo_csv_dumper_52;
    csv_file_dump cstatus_csv_dumper_52;
    df_fifo_monitor fifo_monitor_52;
    df_fifo_intf fifo_intf_53(clock,reset);
    assign fifo_intf_53.rd_en = AESL_inst_myproject.layer4_out_V_2_U.if_read & AESL_inst_myproject.layer4_out_V_2_U.if_empty_n;
    assign fifo_intf_53.wr_en = AESL_inst_myproject.layer4_out_V_2_U.if_write & AESL_inst_myproject.layer4_out_V_2_U.if_full_n;
    assign fifo_intf_53.fifo_rd_block = 0;
    assign fifo_intf_53.fifo_wr_block = 0;
    assign fifo_intf_53.finish = finish;
    csv_file_dump fifo_csv_dumper_53;
    csv_file_dump cstatus_csv_dumper_53;
    df_fifo_monitor fifo_monitor_53;
    df_fifo_intf fifo_intf_54(clock,reset);
    assign fifo_intf_54.rd_en = AESL_inst_myproject.layer4_out_V_3_U.if_read & AESL_inst_myproject.layer4_out_V_3_U.if_empty_n;
    assign fifo_intf_54.wr_en = AESL_inst_myproject.layer4_out_V_3_U.if_write & AESL_inst_myproject.layer4_out_V_3_U.if_full_n;
    assign fifo_intf_54.fifo_rd_block = 0;
    assign fifo_intf_54.fifo_wr_block = 0;
    assign fifo_intf_54.finish = finish;
    csv_file_dump fifo_csv_dumper_54;
    csv_file_dump cstatus_csv_dumper_54;
    df_fifo_monitor fifo_monitor_54;
    df_fifo_intf fifo_intf_55(clock,reset);
    assign fifo_intf_55.rd_en = AESL_inst_myproject.layer4_out_V_4_U.if_read & AESL_inst_myproject.layer4_out_V_4_U.if_empty_n;
    assign fifo_intf_55.wr_en = AESL_inst_myproject.layer4_out_V_4_U.if_write & AESL_inst_myproject.layer4_out_V_4_U.if_full_n;
    assign fifo_intf_55.fifo_rd_block = 0;
    assign fifo_intf_55.fifo_wr_block = 0;
    assign fifo_intf_55.finish = finish;
    csv_file_dump fifo_csv_dumper_55;
    csv_file_dump cstatus_csv_dumper_55;
    df_fifo_monitor fifo_monitor_55;
    df_fifo_intf fifo_intf_56(clock,reset);
    assign fifo_intf_56.rd_en = AESL_inst_myproject.layer4_out_V_5_U.if_read & AESL_inst_myproject.layer4_out_V_5_U.if_empty_n;
    assign fifo_intf_56.wr_en = AESL_inst_myproject.layer4_out_V_5_U.if_write & AESL_inst_myproject.layer4_out_V_5_U.if_full_n;
    assign fifo_intf_56.fifo_rd_block = 0;
    assign fifo_intf_56.fifo_wr_block = 0;
    assign fifo_intf_56.finish = finish;
    csv_file_dump fifo_csv_dumper_56;
    csv_file_dump cstatus_csv_dumper_56;
    df_fifo_monitor fifo_monitor_56;
    df_fifo_intf fifo_intf_57(clock,reset);
    assign fifo_intf_57.rd_en = AESL_inst_myproject.layer4_out_V_6_U.if_read & AESL_inst_myproject.layer4_out_V_6_U.if_empty_n;
    assign fifo_intf_57.wr_en = AESL_inst_myproject.layer4_out_V_6_U.if_write & AESL_inst_myproject.layer4_out_V_6_U.if_full_n;
    assign fifo_intf_57.fifo_rd_block = 0;
    assign fifo_intf_57.fifo_wr_block = 0;
    assign fifo_intf_57.finish = finish;
    csv_file_dump fifo_csv_dumper_57;
    csv_file_dump cstatus_csv_dumper_57;
    df_fifo_monitor fifo_monitor_57;
    df_fifo_intf fifo_intf_58(clock,reset);
    assign fifo_intf_58.rd_en = AESL_inst_myproject.layer4_out_V_7_U.if_read & AESL_inst_myproject.layer4_out_V_7_U.if_empty_n;
    assign fifo_intf_58.wr_en = AESL_inst_myproject.layer4_out_V_7_U.if_write & AESL_inst_myproject.layer4_out_V_7_U.if_full_n;
    assign fifo_intf_58.fifo_rd_block = 0;
    assign fifo_intf_58.fifo_wr_block = 0;
    assign fifo_intf_58.finish = finish;
    csv_file_dump fifo_csv_dumper_58;
    csv_file_dump cstatus_csv_dumper_58;
    df_fifo_monitor fifo_monitor_58;
    df_fifo_intf fifo_intf_59(clock,reset);
    assign fifo_intf_59.rd_en = AESL_inst_myproject.layer4_out_V_8_U.if_read & AESL_inst_myproject.layer4_out_V_8_U.if_empty_n;
    assign fifo_intf_59.wr_en = AESL_inst_myproject.layer4_out_V_8_U.if_write & AESL_inst_myproject.layer4_out_V_8_U.if_full_n;
    assign fifo_intf_59.fifo_rd_block = 0;
    assign fifo_intf_59.fifo_wr_block = 0;
    assign fifo_intf_59.finish = finish;
    csv_file_dump fifo_csv_dumper_59;
    csv_file_dump cstatus_csv_dumper_59;
    df_fifo_monitor fifo_monitor_59;
    df_fifo_intf fifo_intf_60(clock,reset);
    assign fifo_intf_60.rd_en = AESL_inst_myproject.layer4_out_V_9_U.if_read & AESL_inst_myproject.layer4_out_V_9_U.if_empty_n;
    assign fifo_intf_60.wr_en = AESL_inst_myproject.layer4_out_V_9_U.if_write & AESL_inst_myproject.layer4_out_V_9_U.if_full_n;
    assign fifo_intf_60.fifo_rd_block = 0;
    assign fifo_intf_60.fifo_wr_block = 0;
    assign fifo_intf_60.finish = finish;
    csv_file_dump fifo_csv_dumper_60;
    csv_file_dump cstatus_csv_dumper_60;
    df_fifo_monitor fifo_monitor_60;
    df_fifo_intf fifo_intf_61(clock,reset);
    assign fifo_intf_61.rd_en = AESL_inst_myproject.layer4_out_V_10_U.if_read & AESL_inst_myproject.layer4_out_V_10_U.if_empty_n;
    assign fifo_intf_61.wr_en = AESL_inst_myproject.layer4_out_V_10_U.if_write & AESL_inst_myproject.layer4_out_V_10_U.if_full_n;
    assign fifo_intf_61.fifo_rd_block = 0;
    assign fifo_intf_61.fifo_wr_block = 0;
    assign fifo_intf_61.finish = finish;
    csv_file_dump fifo_csv_dumper_61;
    csv_file_dump cstatus_csv_dumper_61;
    df_fifo_monitor fifo_monitor_61;
    df_fifo_intf fifo_intf_62(clock,reset);
    assign fifo_intf_62.rd_en = AESL_inst_myproject.layer4_out_V_11_U.if_read & AESL_inst_myproject.layer4_out_V_11_U.if_empty_n;
    assign fifo_intf_62.wr_en = AESL_inst_myproject.layer4_out_V_11_U.if_write & AESL_inst_myproject.layer4_out_V_11_U.if_full_n;
    assign fifo_intf_62.fifo_rd_block = 0;
    assign fifo_intf_62.fifo_wr_block = 0;
    assign fifo_intf_62.finish = finish;
    csv_file_dump fifo_csv_dumper_62;
    csv_file_dump cstatus_csv_dumper_62;
    df_fifo_monitor fifo_monitor_62;
    df_fifo_intf fifo_intf_63(clock,reset);
    assign fifo_intf_63.rd_en = AESL_inst_myproject.layer4_out_V_12_U.if_read & AESL_inst_myproject.layer4_out_V_12_U.if_empty_n;
    assign fifo_intf_63.wr_en = AESL_inst_myproject.layer4_out_V_12_U.if_write & AESL_inst_myproject.layer4_out_V_12_U.if_full_n;
    assign fifo_intf_63.fifo_rd_block = 0;
    assign fifo_intf_63.fifo_wr_block = 0;
    assign fifo_intf_63.finish = finish;
    csv_file_dump fifo_csv_dumper_63;
    csv_file_dump cstatus_csv_dumper_63;
    df_fifo_monitor fifo_monitor_63;
    df_fifo_intf fifo_intf_64(clock,reset);
    assign fifo_intf_64.rd_en = AESL_inst_myproject.layer4_out_V_13_U.if_read & AESL_inst_myproject.layer4_out_V_13_U.if_empty_n;
    assign fifo_intf_64.wr_en = AESL_inst_myproject.layer4_out_V_13_U.if_write & AESL_inst_myproject.layer4_out_V_13_U.if_full_n;
    assign fifo_intf_64.fifo_rd_block = 0;
    assign fifo_intf_64.fifo_wr_block = 0;
    assign fifo_intf_64.finish = finish;
    csv_file_dump fifo_csv_dumper_64;
    csv_file_dump cstatus_csv_dumper_64;
    df_fifo_monitor fifo_monitor_64;
    df_fifo_intf fifo_intf_65(clock,reset);
    assign fifo_intf_65.rd_en = AESL_inst_myproject.layer4_out_V_14_U.if_read & AESL_inst_myproject.layer4_out_V_14_U.if_empty_n;
    assign fifo_intf_65.wr_en = AESL_inst_myproject.layer4_out_V_14_U.if_write & AESL_inst_myproject.layer4_out_V_14_U.if_full_n;
    assign fifo_intf_65.fifo_rd_block = 0;
    assign fifo_intf_65.fifo_wr_block = 0;
    assign fifo_intf_65.finish = finish;
    csv_file_dump fifo_csv_dumper_65;
    csv_file_dump cstatus_csv_dumper_65;
    df_fifo_monitor fifo_monitor_65;
    df_fifo_intf fifo_intf_66(clock,reset);
    assign fifo_intf_66.rd_en = AESL_inst_myproject.layer4_out_V_15_U.if_read & AESL_inst_myproject.layer4_out_V_15_U.if_empty_n;
    assign fifo_intf_66.wr_en = AESL_inst_myproject.layer4_out_V_15_U.if_write & AESL_inst_myproject.layer4_out_V_15_U.if_full_n;
    assign fifo_intf_66.fifo_rd_block = 0;
    assign fifo_intf_66.fifo_wr_block = 0;
    assign fifo_intf_66.finish = finish;
    csv_file_dump fifo_csv_dumper_66;
    csv_file_dump cstatus_csv_dumper_66;
    df_fifo_monitor fifo_monitor_66;
    df_fifo_intf fifo_intf_67(clock,reset);
    assign fifo_intf_67.rd_en = AESL_inst_myproject.layer4_out_V_16_U.if_read & AESL_inst_myproject.layer4_out_V_16_U.if_empty_n;
    assign fifo_intf_67.wr_en = AESL_inst_myproject.layer4_out_V_16_U.if_write & AESL_inst_myproject.layer4_out_V_16_U.if_full_n;
    assign fifo_intf_67.fifo_rd_block = 0;
    assign fifo_intf_67.fifo_wr_block = 0;
    assign fifo_intf_67.finish = finish;
    csv_file_dump fifo_csv_dumper_67;
    csv_file_dump cstatus_csv_dumper_67;
    df_fifo_monitor fifo_monitor_67;
    df_fifo_intf fifo_intf_68(clock,reset);
    assign fifo_intf_68.rd_en = AESL_inst_myproject.layer4_out_V_17_U.if_read & AESL_inst_myproject.layer4_out_V_17_U.if_empty_n;
    assign fifo_intf_68.wr_en = AESL_inst_myproject.layer4_out_V_17_U.if_write & AESL_inst_myproject.layer4_out_V_17_U.if_full_n;
    assign fifo_intf_68.fifo_rd_block = 0;
    assign fifo_intf_68.fifo_wr_block = 0;
    assign fifo_intf_68.finish = finish;
    csv_file_dump fifo_csv_dumper_68;
    csv_file_dump cstatus_csv_dumper_68;
    df_fifo_monitor fifo_monitor_68;
    df_fifo_intf fifo_intf_69(clock,reset);
    assign fifo_intf_69.rd_en = AESL_inst_myproject.layer4_out_V_18_U.if_read & AESL_inst_myproject.layer4_out_V_18_U.if_empty_n;
    assign fifo_intf_69.wr_en = AESL_inst_myproject.layer4_out_V_18_U.if_write & AESL_inst_myproject.layer4_out_V_18_U.if_full_n;
    assign fifo_intf_69.fifo_rd_block = 0;
    assign fifo_intf_69.fifo_wr_block = 0;
    assign fifo_intf_69.finish = finish;
    csv_file_dump fifo_csv_dumper_69;
    csv_file_dump cstatus_csv_dumper_69;
    df_fifo_monitor fifo_monitor_69;
    df_fifo_intf fifo_intf_70(clock,reset);
    assign fifo_intf_70.rd_en = AESL_inst_myproject.layer4_out_V_19_U.if_read & AESL_inst_myproject.layer4_out_V_19_U.if_empty_n;
    assign fifo_intf_70.wr_en = AESL_inst_myproject.layer4_out_V_19_U.if_write & AESL_inst_myproject.layer4_out_V_19_U.if_full_n;
    assign fifo_intf_70.fifo_rd_block = 0;
    assign fifo_intf_70.fifo_wr_block = 0;
    assign fifo_intf_70.finish = finish;
    csv_file_dump fifo_csv_dumper_70;
    csv_file_dump cstatus_csv_dumper_70;
    df_fifo_monitor fifo_monitor_70;
    df_fifo_intf fifo_intf_71(clock,reset);
    assign fifo_intf_71.rd_en = AESL_inst_myproject.layer4_out_V_20_U.if_read & AESL_inst_myproject.layer4_out_V_20_U.if_empty_n;
    assign fifo_intf_71.wr_en = AESL_inst_myproject.layer4_out_V_20_U.if_write & AESL_inst_myproject.layer4_out_V_20_U.if_full_n;
    assign fifo_intf_71.fifo_rd_block = 0;
    assign fifo_intf_71.fifo_wr_block = 0;
    assign fifo_intf_71.finish = finish;
    csv_file_dump fifo_csv_dumper_71;
    csv_file_dump cstatus_csv_dumper_71;
    df_fifo_monitor fifo_monitor_71;
    df_fifo_intf fifo_intf_72(clock,reset);
    assign fifo_intf_72.rd_en = AESL_inst_myproject.layer4_out_V_21_U.if_read & AESL_inst_myproject.layer4_out_V_21_U.if_empty_n;
    assign fifo_intf_72.wr_en = AESL_inst_myproject.layer4_out_V_21_U.if_write & AESL_inst_myproject.layer4_out_V_21_U.if_full_n;
    assign fifo_intf_72.fifo_rd_block = 0;
    assign fifo_intf_72.fifo_wr_block = 0;
    assign fifo_intf_72.finish = finish;
    csv_file_dump fifo_csv_dumper_72;
    csv_file_dump cstatus_csv_dumper_72;
    df_fifo_monitor fifo_monitor_72;
    df_fifo_intf fifo_intf_73(clock,reset);
    assign fifo_intf_73.rd_en = AESL_inst_myproject.layer4_out_V_22_U.if_read & AESL_inst_myproject.layer4_out_V_22_U.if_empty_n;
    assign fifo_intf_73.wr_en = AESL_inst_myproject.layer4_out_V_22_U.if_write & AESL_inst_myproject.layer4_out_V_22_U.if_full_n;
    assign fifo_intf_73.fifo_rd_block = 0;
    assign fifo_intf_73.fifo_wr_block = 0;
    assign fifo_intf_73.finish = finish;
    csv_file_dump fifo_csv_dumper_73;
    csv_file_dump cstatus_csv_dumper_73;
    df_fifo_monitor fifo_monitor_73;
    df_fifo_intf fifo_intf_74(clock,reset);
    assign fifo_intf_74.rd_en = AESL_inst_myproject.layer4_out_V_23_U.if_read & AESL_inst_myproject.layer4_out_V_23_U.if_empty_n;
    assign fifo_intf_74.wr_en = AESL_inst_myproject.layer4_out_V_23_U.if_write & AESL_inst_myproject.layer4_out_V_23_U.if_full_n;
    assign fifo_intf_74.fifo_rd_block = 0;
    assign fifo_intf_74.fifo_wr_block = 0;
    assign fifo_intf_74.finish = finish;
    csv_file_dump fifo_csv_dumper_74;
    csv_file_dump cstatus_csv_dumper_74;
    df_fifo_monitor fifo_monitor_74;
    df_fifo_intf fifo_intf_75(clock,reset);
    assign fifo_intf_75.rd_en = AESL_inst_myproject.layer4_out_V_24_U.if_read & AESL_inst_myproject.layer4_out_V_24_U.if_empty_n;
    assign fifo_intf_75.wr_en = AESL_inst_myproject.layer4_out_V_24_U.if_write & AESL_inst_myproject.layer4_out_V_24_U.if_full_n;
    assign fifo_intf_75.fifo_rd_block = 0;
    assign fifo_intf_75.fifo_wr_block = 0;
    assign fifo_intf_75.finish = finish;
    csv_file_dump fifo_csv_dumper_75;
    csv_file_dump cstatus_csv_dumper_75;
    df_fifo_monitor fifo_monitor_75;
    df_fifo_intf fifo_intf_76(clock,reset);
    assign fifo_intf_76.rd_en = AESL_inst_myproject.layer4_out_V_25_U.if_read & AESL_inst_myproject.layer4_out_V_25_U.if_empty_n;
    assign fifo_intf_76.wr_en = AESL_inst_myproject.layer4_out_V_25_U.if_write & AESL_inst_myproject.layer4_out_V_25_U.if_full_n;
    assign fifo_intf_76.fifo_rd_block = 0;
    assign fifo_intf_76.fifo_wr_block = 0;
    assign fifo_intf_76.finish = finish;
    csv_file_dump fifo_csv_dumper_76;
    csv_file_dump cstatus_csv_dumper_76;
    df_fifo_monitor fifo_monitor_76;
    df_fifo_intf fifo_intf_77(clock,reset);
    assign fifo_intf_77.rd_en = AESL_inst_myproject.layer4_out_V_26_U.if_read & AESL_inst_myproject.layer4_out_V_26_U.if_empty_n;
    assign fifo_intf_77.wr_en = AESL_inst_myproject.layer4_out_V_26_U.if_write & AESL_inst_myproject.layer4_out_V_26_U.if_full_n;
    assign fifo_intf_77.fifo_rd_block = 0;
    assign fifo_intf_77.fifo_wr_block = 0;
    assign fifo_intf_77.finish = finish;
    csv_file_dump fifo_csv_dumper_77;
    csv_file_dump cstatus_csv_dumper_77;
    df_fifo_monitor fifo_monitor_77;
    df_fifo_intf fifo_intf_78(clock,reset);
    assign fifo_intf_78.rd_en = AESL_inst_myproject.layer4_out_V_27_U.if_read & AESL_inst_myproject.layer4_out_V_27_U.if_empty_n;
    assign fifo_intf_78.wr_en = AESL_inst_myproject.layer4_out_V_27_U.if_write & AESL_inst_myproject.layer4_out_V_27_U.if_full_n;
    assign fifo_intf_78.fifo_rd_block = 0;
    assign fifo_intf_78.fifo_wr_block = 0;
    assign fifo_intf_78.finish = finish;
    csv_file_dump fifo_csv_dumper_78;
    csv_file_dump cstatus_csv_dumper_78;
    df_fifo_monitor fifo_monitor_78;
    df_fifo_intf fifo_intf_79(clock,reset);
    assign fifo_intf_79.rd_en = AESL_inst_myproject.layer4_out_V_28_U.if_read & AESL_inst_myproject.layer4_out_V_28_U.if_empty_n;
    assign fifo_intf_79.wr_en = AESL_inst_myproject.layer4_out_V_28_U.if_write & AESL_inst_myproject.layer4_out_V_28_U.if_full_n;
    assign fifo_intf_79.fifo_rd_block = 0;
    assign fifo_intf_79.fifo_wr_block = 0;
    assign fifo_intf_79.finish = finish;
    csv_file_dump fifo_csv_dumper_79;
    csv_file_dump cstatus_csv_dumper_79;
    df_fifo_monitor fifo_monitor_79;
    df_fifo_intf fifo_intf_80(clock,reset);
    assign fifo_intf_80.rd_en = AESL_inst_myproject.layer4_out_V_29_U.if_read & AESL_inst_myproject.layer4_out_V_29_U.if_empty_n;
    assign fifo_intf_80.wr_en = AESL_inst_myproject.layer4_out_V_29_U.if_write & AESL_inst_myproject.layer4_out_V_29_U.if_full_n;
    assign fifo_intf_80.fifo_rd_block = 0;
    assign fifo_intf_80.fifo_wr_block = 0;
    assign fifo_intf_80.finish = finish;
    csv_file_dump fifo_csv_dumper_80;
    csv_file_dump cstatus_csv_dumper_80;
    df_fifo_monitor fifo_monitor_80;
    df_fifo_intf fifo_intf_81(clock,reset);
    assign fifo_intf_81.rd_en = AESL_inst_myproject.layer4_out_V_30_U.if_read & AESL_inst_myproject.layer4_out_V_30_U.if_empty_n;
    assign fifo_intf_81.wr_en = AESL_inst_myproject.layer4_out_V_30_U.if_write & AESL_inst_myproject.layer4_out_V_30_U.if_full_n;
    assign fifo_intf_81.fifo_rd_block = 0;
    assign fifo_intf_81.fifo_wr_block = 0;
    assign fifo_intf_81.finish = finish;
    csv_file_dump fifo_csv_dumper_81;
    csv_file_dump cstatus_csv_dumper_81;
    df_fifo_monitor fifo_monitor_81;
    df_fifo_intf fifo_intf_82(clock,reset);
    assign fifo_intf_82.rd_en = AESL_inst_myproject.layer4_out_V_31_U.if_read & AESL_inst_myproject.layer4_out_V_31_U.if_empty_n;
    assign fifo_intf_82.wr_en = AESL_inst_myproject.layer4_out_V_31_U.if_write & AESL_inst_myproject.layer4_out_V_31_U.if_full_n;
    assign fifo_intf_82.fifo_rd_block = 0;
    assign fifo_intf_82.fifo_wr_block = 0;
    assign fifo_intf_82.finish = finish;
    csv_file_dump fifo_csv_dumper_82;
    csv_file_dump cstatus_csv_dumper_82;
    df_fifo_monitor fifo_monitor_82;
    df_fifo_intf fifo_intf_83(clock,reset);
    assign fifo_intf_83.rd_en = AESL_inst_myproject.layer4_out_V_32_U.if_read & AESL_inst_myproject.layer4_out_V_32_U.if_empty_n;
    assign fifo_intf_83.wr_en = AESL_inst_myproject.layer4_out_V_32_U.if_write & AESL_inst_myproject.layer4_out_V_32_U.if_full_n;
    assign fifo_intf_83.fifo_rd_block = 0;
    assign fifo_intf_83.fifo_wr_block = 0;
    assign fifo_intf_83.finish = finish;
    csv_file_dump fifo_csv_dumper_83;
    csv_file_dump cstatus_csv_dumper_83;
    df_fifo_monitor fifo_monitor_83;
    df_fifo_intf fifo_intf_84(clock,reset);
    assign fifo_intf_84.rd_en = AESL_inst_myproject.layer4_out_V_33_U.if_read & AESL_inst_myproject.layer4_out_V_33_U.if_empty_n;
    assign fifo_intf_84.wr_en = AESL_inst_myproject.layer4_out_V_33_U.if_write & AESL_inst_myproject.layer4_out_V_33_U.if_full_n;
    assign fifo_intf_84.fifo_rd_block = 0;
    assign fifo_intf_84.fifo_wr_block = 0;
    assign fifo_intf_84.finish = finish;
    csv_file_dump fifo_csv_dumper_84;
    csv_file_dump cstatus_csv_dumper_84;
    df_fifo_monitor fifo_monitor_84;
    df_fifo_intf fifo_intf_85(clock,reset);
    assign fifo_intf_85.rd_en = AESL_inst_myproject.layer4_out_V_34_U.if_read & AESL_inst_myproject.layer4_out_V_34_U.if_empty_n;
    assign fifo_intf_85.wr_en = AESL_inst_myproject.layer4_out_V_34_U.if_write & AESL_inst_myproject.layer4_out_V_34_U.if_full_n;
    assign fifo_intf_85.fifo_rd_block = 0;
    assign fifo_intf_85.fifo_wr_block = 0;
    assign fifo_intf_85.finish = finish;
    csv_file_dump fifo_csv_dumper_85;
    csv_file_dump cstatus_csv_dumper_85;
    df_fifo_monitor fifo_monitor_85;
    df_fifo_intf fifo_intf_86(clock,reset);
    assign fifo_intf_86.rd_en = AESL_inst_myproject.layer4_out_V_35_U.if_read & AESL_inst_myproject.layer4_out_V_35_U.if_empty_n;
    assign fifo_intf_86.wr_en = AESL_inst_myproject.layer4_out_V_35_U.if_write & AESL_inst_myproject.layer4_out_V_35_U.if_full_n;
    assign fifo_intf_86.fifo_rd_block = 0;
    assign fifo_intf_86.fifo_wr_block = 0;
    assign fifo_intf_86.finish = finish;
    csv_file_dump fifo_csv_dumper_86;
    csv_file_dump cstatus_csv_dumper_86;
    df_fifo_monitor fifo_monitor_86;
    df_fifo_intf fifo_intf_87(clock,reset);
    assign fifo_intf_87.rd_en = AESL_inst_myproject.layer4_out_V_36_U.if_read & AESL_inst_myproject.layer4_out_V_36_U.if_empty_n;
    assign fifo_intf_87.wr_en = AESL_inst_myproject.layer4_out_V_36_U.if_write & AESL_inst_myproject.layer4_out_V_36_U.if_full_n;
    assign fifo_intf_87.fifo_rd_block = 0;
    assign fifo_intf_87.fifo_wr_block = 0;
    assign fifo_intf_87.finish = finish;
    csv_file_dump fifo_csv_dumper_87;
    csv_file_dump cstatus_csv_dumper_87;
    df_fifo_monitor fifo_monitor_87;
    df_fifo_intf fifo_intf_88(clock,reset);
    assign fifo_intf_88.rd_en = AESL_inst_myproject.layer4_out_V_37_U.if_read & AESL_inst_myproject.layer4_out_V_37_U.if_empty_n;
    assign fifo_intf_88.wr_en = AESL_inst_myproject.layer4_out_V_37_U.if_write & AESL_inst_myproject.layer4_out_V_37_U.if_full_n;
    assign fifo_intf_88.fifo_rd_block = 0;
    assign fifo_intf_88.fifo_wr_block = 0;
    assign fifo_intf_88.finish = finish;
    csv_file_dump fifo_csv_dumper_88;
    csv_file_dump cstatus_csv_dumper_88;
    df_fifo_monitor fifo_monitor_88;
    df_fifo_intf fifo_intf_89(clock,reset);
    assign fifo_intf_89.rd_en = AESL_inst_myproject.layer4_out_V_38_U.if_read & AESL_inst_myproject.layer4_out_V_38_U.if_empty_n;
    assign fifo_intf_89.wr_en = AESL_inst_myproject.layer4_out_V_38_U.if_write & AESL_inst_myproject.layer4_out_V_38_U.if_full_n;
    assign fifo_intf_89.fifo_rd_block = 0;
    assign fifo_intf_89.fifo_wr_block = 0;
    assign fifo_intf_89.finish = finish;
    csv_file_dump fifo_csv_dumper_89;
    csv_file_dump cstatus_csv_dumper_89;
    df_fifo_monitor fifo_monitor_89;
    df_fifo_intf fifo_intf_90(clock,reset);
    assign fifo_intf_90.rd_en = AESL_inst_myproject.layer4_out_V_39_U.if_read & AESL_inst_myproject.layer4_out_V_39_U.if_empty_n;
    assign fifo_intf_90.wr_en = AESL_inst_myproject.layer4_out_V_39_U.if_write & AESL_inst_myproject.layer4_out_V_39_U.if_full_n;
    assign fifo_intf_90.fifo_rd_block = 0;
    assign fifo_intf_90.fifo_wr_block = 0;
    assign fifo_intf_90.finish = finish;
    csv_file_dump fifo_csv_dumper_90;
    csv_file_dump cstatus_csv_dumper_90;
    df_fifo_monitor fifo_monitor_90;
    df_fifo_intf fifo_intf_91(clock,reset);
    assign fifo_intf_91.rd_en = AESL_inst_myproject.layer4_out_V_40_U.if_read & AESL_inst_myproject.layer4_out_V_40_U.if_empty_n;
    assign fifo_intf_91.wr_en = AESL_inst_myproject.layer4_out_V_40_U.if_write & AESL_inst_myproject.layer4_out_V_40_U.if_full_n;
    assign fifo_intf_91.fifo_rd_block = 0;
    assign fifo_intf_91.fifo_wr_block = 0;
    assign fifo_intf_91.finish = finish;
    csv_file_dump fifo_csv_dumper_91;
    csv_file_dump cstatus_csv_dumper_91;
    df_fifo_monitor fifo_monitor_91;
    df_fifo_intf fifo_intf_92(clock,reset);
    assign fifo_intf_92.rd_en = AESL_inst_myproject.layer4_out_V_41_U.if_read & AESL_inst_myproject.layer4_out_V_41_U.if_empty_n;
    assign fifo_intf_92.wr_en = AESL_inst_myproject.layer4_out_V_41_U.if_write & AESL_inst_myproject.layer4_out_V_41_U.if_full_n;
    assign fifo_intf_92.fifo_rd_block = 0;
    assign fifo_intf_92.fifo_wr_block = 0;
    assign fifo_intf_92.finish = finish;
    csv_file_dump fifo_csv_dumper_92;
    csv_file_dump cstatus_csv_dumper_92;
    df_fifo_monitor fifo_monitor_92;
    df_fifo_intf fifo_intf_93(clock,reset);
    assign fifo_intf_93.rd_en = AESL_inst_myproject.layer4_out_V_42_U.if_read & AESL_inst_myproject.layer4_out_V_42_U.if_empty_n;
    assign fifo_intf_93.wr_en = AESL_inst_myproject.layer4_out_V_42_U.if_write & AESL_inst_myproject.layer4_out_V_42_U.if_full_n;
    assign fifo_intf_93.fifo_rd_block = 0;
    assign fifo_intf_93.fifo_wr_block = 0;
    assign fifo_intf_93.finish = finish;
    csv_file_dump fifo_csv_dumper_93;
    csv_file_dump cstatus_csv_dumper_93;
    df_fifo_monitor fifo_monitor_93;
    df_fifo_intf fifo_intf_94(clock,reset);
    assign fifo_intf_94.rd_en = AESL_inst_myproject.layer4_out_V_43_U.if_read & AESL_inst_myproject.layer4_out_V_43_U.if_empty_n;
    assign fifo_intf_94.wr_en = AESL_inst_myproject.layer4_out_V_43_U.if_write & AESL_inst_myproject.layer4_out_V_43_U.if_full_n;
    assign fifo_intf_94.fifo_rd_block = 0;
    assign fifo_intf_94.fifo_wr_block = 0;
    assign fifo_intf_94.finish = finish;
    csv_file_dump fifo_csv_dumper_94;
    csv_file_dump cstatus_csv_dumper_94;
    df_fifo_monitor fifo_monitor_94;
    df_fifo_intf fifo_intf_95(clock,reset);
    assign fifo_intf_95.rd_en = AESL_inst_myproject.layer4_out_V_44_U.if_read & AESL_inst_myproject.layer4_out_V_44_U.if_empty_n;
    assign fifo_intf_95.wr_en = AESL_inst_myproject.layer4_out_V_44_U.if_write & AESL_inst_myproject.layer4_out_V_44_U.if_full_n;
    assign fifo_intf_95.fifo_rd_block = 0;
    assign fifo_intf_95.fifo_wr_block = 0;
    assign fifo_intf_95.finish = finish;
    csv_file_dump fifo_csv_dumper_95;
    csv_file_dump cstatus_csv_dumper_95;
    df_fifo_monitor fifo_monitor_95;
    df_fifo_intf fifo_intf_96(clock,reset);
    assign fifo_intf_96.rd_en = AESL_inst_myproject.layer4_out_V_45_U.if_read & AESL_inst_myproject.layer4_out_V_45_U.if_empty_n;
    assign fifo_intf_96.wr_en = AESL_inst_myproject.layer4_out_V_45_U.if_write & AESL_inst_myproject.layer4_out_V_45_U.if_full_n;
    assign fifo_intf_96.fifo_rd_block = 0;
    assign fifo_intf_96.fifo_wr_block = 0;
    assign fifo_intf_96.finish = finish;
    csv_file_dump fifo_csv_dumper_96;
    csv_file_dump cstatus_csv_dumper_96;
    df_fifo_monitor fifo_monitor_96;
    df_fifo_intf fifo_intf_97(clock,reset);
    assign fifo_intf_97.rd_en = AESL_inst_myproject.layer4_out_V_46_U.if_read & AESL_inst_myproject.layer4_out_V_46_U.if_empty_n;
    assign fifo_intf_97.wr_en = AESL_inst_myproject.layer4_out_V_46_U.if_write & AESL_inst_myproject.layer4_out_V_46_U.if_full_n;
    assign fifo_intf_97.fifo_rd_block = 0;
    assign fifo_intf_97.fifo_wr_block = 0;
    assign fifo_intf_97.finish = finish;
    csv_file_dump fifo_csv_dumper_97;
    csv_file_dump cstatus_csv_dumper_97;
    df_fifo_monitor fifo_monitor_97;
    df_fifo_intf fifo_intf_98(clock,reset);
    assign fifo_intf_98.rd_en = AESL_inst_myproject.layer4_out_V_47_U.if_read & AESL_inst_myproject.layer4_out_V_47_U.if_empty_n;
    assign fifo_intf_98.wr_en = AESL_inst_myproject.layer4_out_V_47_U.if_write & AESL_inst_myproject.layer4_out_V_47_U.if_full_n;
    assign fifo_intf_98.fifo_rd_block = 0;
    assign fifo_intf_98.fifo_wr_block = 0;
    assign fifo_intf_98.finish = finish;
    csv_file_dump fifo_csv_dumper_98;
    csv_file_dump cstatus_csv_dumper_98;
    df_fifo_monitor fifo_monitor_98;
    df_fifo_intf fifo_intf_99(clock,reset);
    assign fifo_intf_99.rd_en = AESL_inst_myproject.layer4_out_V_48_U.if_read & AESL_inst_myproject.layer4_out_V_48_U.if_empty_n;
    assign fifo_intf_99.wr_en = AESL_inst_myproject.layer4_out_V_48_U.if_write & AESL_inst_myproject.layer4_out_V_48_U.if_full_n;
    assign fifo_intf_99.fifo_rd_block = 0;
    assign fifo_intf_99.fifo_wr_block = 0;
    assign fifo_intf_99.finish = finish;
    csv_file_dump fifo_csv_dumper_99;
    csv_file_dump cstatus_csv_dumper_99;
    df_fifo_monitor fifo_monitor_99;
    df_fifo_intf fifo_intf_100(clock,reset);
    assign fifo_intf_100.rd_en = AESL_inst_myproject.layer4_out_V_49_U.if_read & AESL_inst_myproject.layer4_out_V_49_U.if_empty_n;
    assign fifo_intf_100.wr_en = AESL_inst_myproject.layer4_out_V_49_U.if_write & AESL_inst_myproject.layer4_out_V_49_U.if_full_n;
    assign fifo_intf_100.fifo_rd_block = 0;
    assign fifo_intf_100.fifo_wr_block = 0;
    assign fifo_intf_100.finish = finish;
    csv_file_dump fifo_csv_dumper_100;
    csv_file_dump cstatus_csv_dumper_100;
    df_fifo_monitor fifo_monitor_100;
    df_fifo_intf fifo_intf_101(clock,reset);
    assign fifo_intf_101.rd_en = AESL_inst_myproject.layer5_out_V_U.if_read & AESL_inst_myproject.layer5_out_V_U.if_empty_n;
    assign fifo_intf_101.wr_en = AESL_inst_myproject.layer5_out_V_U.if_write & AESL_inst_myproject.layer5_out_V_U.if_full_n;
    assign fifo_intf_101.fifo_rd_block = 0;
    assign fifo_intf_101.fifo_wr_block = 0;
    assign fifo_intf_101.finish = finish;
    csv_file_dump fifo_csv_dumper_101;
    csv_file_dump cstatus_csv_dumper_101;
    df_fifo_monitor fifo_monitor_101;
    df_fifo_intf fifo_intf_102(clock,reset);
    assign fifo_intf_102.rd_en = AESL_inst_myproject.layer5_out_V_1_U.if_read & AESL_inst_myproject.layer5_out_V_1_U.if_empty_n;
    assign fifo_intf_102.wr_en = AESL_inst_myproject.layer5_out_V_1_U.if_write & AESL_inst_myproject.layer5_out_V_1_U.if_full_n;
    assign fifo_intf_102.fifo_rd_block = 0;
    assign fifo_intf_102.fifo_wr_block = 0;
    assign fifo_intf_102.finish = finish;
    csv_file_dump fifo_csv_dumper_102;
    csv_file_dump cstatus_csv_dumper_102;
    df_fifo_monitor fifo_monitor_102;
    df_fifo_intf fifo_intf_103(clock,reset);
    assign fifo_intf_103.rd_en = AESL_inst_myproject.layer5_out_V_2_U.if_read & AESL_inst_myproject.layer5_out_V_2_U.if_empty_n;
    assign fifo_intf_103.wr_en = AESL_inst_myproject.layer5_out_V_2_U.if_write & AESL_inst_myproject.layer5_out_V_2_U.if_full_n;
    assign fifo_intf_103.fifo_rd_block = 0;
    assign fifo_intf_103.fifo_wr_block = 0;
    assign fifo_intf_103.finish = finish;
    csv_file_dump fifo_csv_dumper_103;
    csv_file_dump cstatus_csv_dumper_103;
    df_fifo_monitor fifo_monitor_103;
    df_fifo_intf fifo_intf_104(clock,reset);
    assign fifo_intf_104.rd_en = AESL_inst_myproject.layer5_out_V_3_U.if_read & AESL_inst_myproject.layer5_out_V_3_U.if_empty_n;
    assign fifo_intf_104.wr_en = AESL_inst_myproject.layer5_out_V_3_U.if_write & AESL_inst_myproject.layer5_out_V_3_U.if_full_n;
    assign fifo_intf_104.fifo_rd_block = 0;
    assign fifo_intf_104.fifo_wr_block = 0;
    assign fifo_intf_104.finish = finish;
    csv_file_dump fifo_csv_dumper_104;
    csv_file_dump cstatus_csv_dumper_104;
    df_fifo_monitor fifo_monitor_104;
    df_fifo_intf fifo_intf_105(clock,reset);
    assign fifo_intf_105.rd_en = AESL_inst_myproject.layer5_out_V_4_U.if_read & AESL_inst_myproject.layer5_out_V_4_U.if_empty_n;
    assign fifo_intf_105.wr_en = AESL_inst_myproject.layer5_out_V_4_U.if_write & AESL_inst_myproject.layer5_out_V_4_U.if_full_n;
    assign fifo_intf_105.fifo_rd_block = 0;
    assign fifo_intf_105.fifo_wr_block = 0;
    assign fifo_intf_105.finish = finish;
    csv_file_dump fifo_csv_dumper_105;
    csv_file_dump cstatus_csv_dumper_105;
    df_fifo_monitor fifo_monitor_105;
    df_fifo_intf fifo_intf_106(clock,reset);
    assign fifo_intf_106.rd_en = AESL_inst_myproject.layer5_out_V_5_U.if_read & AESL_inst_myproject.layer5_out_V_5_U.if_empty_n;
    assign fifo_intf_106.wr_en = AESL_inst_myproject.layer5_out_V_5_U.if_write & AESL_inst_myproject.layer5_out_V_5_U.if_full_n;
    assign fifo_intf_106.fifo_rd_block = 0;
    assign fifo_intf_106.fifo_wr_block = 0;
    assign fifo_intf_106.finish = finish;
    csv_file_dump fifo_csv_dumper_106;
    csv_file_dump cstatus_csv_dumper_106;
    df_fifo_monitor fifo_monitor_106;
    df_fifo_intf fifo_intf_107(clock,reset);
    assign fifo_intf_107.rd_en = AESL_inst_myproject.layer5_out_V_6_U.if_read & AESL_inst_myproject.layer5_out_V_6_U.if_empty_n;
    assign fifo_intf_107.wr_en = AESL_inst_myproject.layer5_out_V_6_U.if_write & AESL_inst_myproject.layer5_out_V_6_U.if_full_n;
    assign fifo_intf_107.fifo_rd_block = 0;
    assign fifo_intf_107.fifo_wr_block = 0;
    assign fifo_intf_107.finish = finish;
    csv_file_dump fifo_csv_dumper_107;
    csv_file_dump cstatus_csv_dumper_107;
    df_fifo_monitor fifo_monitor_107;
    df_fifo_intf fifo_intf_108(clock,reset);
    assign fifo_intf_108.rd_en = AESL_inst_myproject.layer5_out_V_7_U.if_read & AESL_inst_myproject.layer5_out_V_7_U.if_empty_n;
    assign fifo_intf_108.wr_en = AESL_inst_myproject.layer5_out_V_7_U.if_write & AESL_inst_myproject.layer5_out_V_7_U.if_full_n;
    assign fifo_intf_108.fifo_rd_block = 0;
    assign fifo_intf_108.fifo_wr_block = 0;
    assign fifo_intf_108.finish = finish;
    csv_file_dump fifo_csv_dumper_108;
    csv_file_dump cstatus_csv_dumper_108;
    df_fifo_monitor fifo_monitor_108;
    df_fifo_intf fifo_intf_109(clock,reset);
    assign fifo_intf_109.rd_en = AESL_inst_myproject.layer5_out_V_8_U.if_read & AESL_inst_myproject.layer5_out_V_8_U.if_empty_n;
    assign fifo_intf_109.wr_en = AESL_inst_myproject.layer5_out_V_8_U.if_write & AESL_inst_myproject.layer5_out_V_8_U.if_full_n;
    assign fifo_intf_109.fifo_rd_block = 0;
    assign fifo_intf_109.fifo_wr_block = 0;
    assign fifo_intf_109.finish = finish;
    csv_file_dump fifo_csv_dumper_109;
    csv_file_dump cstatus_csv_dumper_109;
    df_fifo_monitor fifo_monitor_109;
    df_fifo_intf fifo_intf_110(clock,reset);
    assign fifo_intf_110.rd_en = AESL_inst_myproject.layer5_out_V_9_U.if_read & AESL_inst_myproject.layer5_out_V_9_U.if_empty_n;
    assign fifo_intf_110.wr_en = AESL_inst_myproject.layer5_out_V_9_U.if_write & AESL_inst_myproject.layer5_out_V_9_U.if_full_n;
    assign fifo_intf_110.fifo_rd_block = 0;
    assign fifo_intf_110.fifo_wr_block = 0;
    assign fifo_intf_110.finish = finish;
    csv_file_dump fifo_csv_dumper_110;
    csv_file_dump cstatus_csv_dumper_110;
    df_fifo_monitor fifo_monitor_110;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_myproject.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_myproject.ap_start == 1'b1 && AESL_inst_myproject.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_myproject.ap_done == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_0_idle;
    assign process_intf_1.finish = finish;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_myproject.relu_ap_fixed_ap_fixed_16_8_5_3_0_relu_config4_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_myproject.relu_ap_fixed_ap_fixed_16_8_5_3_0_relu_config4_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_myproject.relu_ap_fixed_ap_fixed_16_8_5_3_0_relu_config4_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_myproject.relu_ap_fixed_ap_fixed_16_8_5_3_0_relu_config4_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_myproject.relu_ap_fixed_ap_fixed_16_8_5_3_0_relu_config4_U0.ap_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0;
    assign process_intf_2.region_idle = region_0_idle;
    assign process_intf_2.finish = finish;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_start;
    assign process_intf_3.pin_stall = 1'b0;
    assign process_intf_3.pout_stall = 1'b0;
    assign process_intf_3.cin_stall = 1'b0;
    assign process_intf_3.cout_stall = 1'b0;
    assign process_intf_3.region_idle = region_0_idle;
    assign process_intf_3.finish = finish;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_myproject.softmax_latency_ap_fixed_ap_fixed_softmax_config7_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_myproject.softmax_latency_ap_fixed_ap_fixed_softmax_config7_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_myproject.softmax_latency_ap_fixed_ap_fixed_softmax_config7_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_myproject.softmax_latency_ap_fixed_ap_fixed_softmax_config7_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_myproject.softmax_latency_ap_fixed_ap_fixed_softmax_config7_U0.ap_start;
    assign process_intf_4.pin_stall = 1'b0;
    assign process_intf_4.pout_stall = 1'b0;
    assign process_intf_4.cin_stall = 1'b0;
    assign process_intf_4.cout_stall = 1'b0;
    assign process_intf_4.region_idle = region_0_idle;
    assign process_intf_4.finish = finish;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_myproject.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_myproject.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_myproject.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;

    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_1.quit_enable = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_1.loop_start = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_done;
    assign upc_loop_intf_1.loop_continue = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config2_U0.ap_continue;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_2.quit_enable = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_2.loop_start = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_done;
    assign upc_loop_intf_2.loop_continue = AESL_inst_myproject.dense_resource_ap_fixed_ap_fixed_16_8_5_3_0_config5_U0.ap_continue;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);
    fifo_csv_dumper_18 = new("./depth18.csv");
    cstatus_csv_dumper_18 = new("./chan_status18.csv");
    fifo_monitor_18 = new(fifo_csv_dumper_18,fifo_intf_18,cstatus_csv_dumper_18);
    fifo_csv_dumper_19 = new("./depth19.csv");
    cstatus_csv_dumper_19 = new("./chan_status19.csv");
    fifo_monitor_19 = new(fifo_csv_dumper_19,fifo_intf_19,cstatus_csv_dumper_19);
    fifo_csv_dumper_20 = new("./depth20.csv");
    cstatus_csv_dumper_20 = new("./chan_status20.csv");
    fifo_monitor_20 = new(fifo_csv_dumper_20,fifo_intf_20,cstatus_csv_dumper_20);
    fifo_csv_dumper_21 = new("./depth21.csv");
    cstatus_csv_dumper_21 = new("./chan_status21.csv");
    fifo_monitor_21 = new(fifo_csv_dumper_21,fifo_intf_21,cstatus_csv_dumper_21);
    fifo_csv_dumper_22 = new("./depth22.csv");
    cstatus_csv_dumper_22 = new("./chan_status22.csv");
    fifo_monitor_22 = new(fifo_csv_dumper_22,fifo_intf_22,cstatus_csv_dumper_22);
    fifo_csv_dumper_23 = new("./depth23.csv");
    cstatus_csv_dumper_23 = new("./chan_status23.csv");
    fifo_monitor_23 = new(fifo_csv_dumper_23,fifo_intf_23,cstatus_csv_dumper_23);
    fifo_csv_dumper_24 = new("./depth24.csv");
    cstatus_csv_dumper_24 = new("./chan_status24.csv");
    fifo_monitor_24 = new(fifo_csv_dumper_24,fifo_intf_24,cstatus_csv_dumper_24);
    fifo_csv_dumper_25 = new("./depth25.csv");
    cstatus_csv_dumper_25 = new("./chan_status25.csv");
    fifo_monitor_25 = new(fifo_csv_dumper_25,fifo_intf_25,cstatus_csv_dumper_25);
    fifo_csv_dumper_26 = new("./depth26.csv");
    cstatus_csv_dumper_26 = new("./chan_status26.csv");
    fifo_monitor_26 = new(fifo_csv_dumper_26,fifo_intf_26,cstatus_csv_dumper_26);
    fifo_csv_dumper_27 = new("./depth27.csv");
    cstatus_csv_dumper_27 = new("./chan_status27.csv");
    fifo_monitor_27 = new(fifo_csv_dumper_27,fifo_intf_27,cstatus_csv_dumper_27);
    fifo_csv_dumper_28 = new("./depth28.csv");
    cstatus_csv_dumper_28 = new("./chan_status28.csv");
    fifo_monitor_28 = new(fifo_csv_dumper_28,fifo_intf_28,cstatus_csv_dumper_28);
    fifo_csv_dumper_29 = new("./depth29.csv");
    cstatus_csv_dumper_29 = new("./chan_status29.csv");
    fifo_monitor_29 = new(fifo_csv_dumper_29,fifo_intf_29,cstatus_csv_dumper_29);
    fifo_csv_dumper_30 = new("./depth30.csv");
    cstatus_csv_dumper_30 = new("./chan_status30.csv");
    fifo_monitor_30 = new(fifo_csv_dumper_30,fifo_intf_30,cstatus_csv_dumper_30);
    fifo_csv_dumper_31 = new("./depth31.csv");
    cstatus_csv_dumper_31 = new("./chan_status31.csv");
    fifo_monitor_31 = new(fifo_csv_dumper_31,fifo_intf_31,cstatus_csv_dumper_31);
    fifo_csv_dumper_32 = new("./depth32.csv");
    cstatus_csv_dumper_32 = new("./chan_status32.csv");
    fifo_monitor_32 = new(fifo_csv_dumper_32,fifo_intf_32,cstatus_csv_dumper_32);
    fifo_csv_dumper_33 = new("./depth33.csv");
    cstatus_csv_dumper_33 = new("./chan_status33.csv");
    fifo_monitor_33 = new(fifo_csv_dumper_33,fifo_intf_33,cstatus_csv_dumper_33);
    fifo_csv_dumper_34 = new("./depth34.csv");
    cstatus_csv_dumper_34 = new("./chan_status34.csv");
    fifo_monitor_34 = new(fifo_csv_dumper_34,fifo_intf_34,cstatus_csv_dumper_34);
    fifo_csv_dumper_35 = new("./depth35.csv");
    cstatus_csv_dumper_35 = new("./chan_status35.csv");
    fifo_monitor_35 = new(fifo_csv_dumper_35,fifo_intf_35,cstatus_csv_dumper_35);
    fifo_csv_dumper_36 = new("./depth36.csv");
    cstatus_csv_dumper_36 = new("./chan_status36.csv");
    fifo_monitor_36 = new(fifo_csv_dumper_36,fifo_intf_36,cstatus_csv_dumper_36);
    fifo_csv_dumper_37 = new("./depth37.csv");
    cstatus_csv_dumper_37 = new("./chan_status37.csv");
    fifo_monitor_37 = new(fifo_csv_dumper_37,fifo_intf_37,cstatus_csv_dumper_37);
    fifo_csv_dumper_38 = new("./depth38.csv");
    cstatus_csv_dumper_38 = new("./chan_status38.csv");
    fifo_monitor_38 = new(fifo_csv_dumper_38,fifo_intf_38,cstatus_csv_dumper_38);
    fifo_csv_dumper_39 = new("./depth39.csv");
    cstatus_csv_dumper_39 = new("./chan_status39.csv");
    fifo_monitor_39 = new(fifo_csv_dumper_39,fifo_intf_39,cstatus_csv_dumper_39);
    fifo_csv_dumper_40 = new("./depth40.csv");
    cstatus_csv_dumper_40 = new("./chan_status40.csv");
    fifo_monitor_40 = new(fifo_csv_dumper_40,fifo_intf_40,cstatus_csv_dumper_40);
    fifo_csv_dumper_41 = new("./depth41.csv");
    cstatus_csv_dumper_41 = new("./chan_status41.csv");
    fifo_monitor_41 = new(fifo_csv_dumper_41,fifo_intf_41,cstatus_csv_dumper_41);
    fifo_csv_dumper_42 = new("./depth42.csv");
    cstatus_csv_dumper_42 = new("./chan_status42.csv");
    fifo_monitor_42 = new(fifo_csv_dumper_42,fifo_intf_42,cstatus_csv_dumper_42);
    fifo_csv_dumper_43 = new("./depth43.csv");
    cstatus_csv_dumper_43 = new("./chan_status43.csv");
    fifo_monitor_43 = new(fifo_csv_dumper_43,fifo_intf_43,cstatus_csv_dumper_43);
    fifo_csv_dumper_44 = new("./depth44.csv");
    cstatus_csv_dumper_44 = new("./chan_status44.csv");
    fifo_monitor_44 = new(fifo_csv_dumper_44,fifo_intf_44,cstatus_csv_dumper_44);
    fifo_csv_dumper_45 = new("./depth45.csv");
    cstatus_csv_dumper_45 = new("./chan_status45.csv");
    fifo_monitor_45 = new(fifo_csv_dumper_45,fifo_intf_45,cstatus_csv_dumper_45);
    fifo_csv_dumper_46 = new("./depth46.csv");
    cstatus_csv_dumper_46 = new("./chan_status46.csv");
    fifo_monitor_46 = new(fifo_csv_dumper_46,fifo_intf_46,cstatus_csv_dumper_46);
    fifo_csv_dumper_47 = new("./depth47.csv");
    cstatus_csv_dumper_47 = new("./chan_status47.csv");
    fifo_monitor_47 = new(fifo_csv_dumper_47,fifo_intf_47,cstatus_csv_dumper_47);
    fifo_csv_dumper_48 = new("./depth48.csv");
    cstatus_csv_dumper_48 = new("./chan_status48.csv");
    fifo_monitor_48 = new(fifo_csv_dumper_48,fifo_intf_48,cstatus_csv_dumper_48);
    fifo_csv_dumper_49 = new("./depth49.csv");
    cstatus_csv_dumper_49 = new("./chan_status49.csv");
    fifo_monitor_49 = new(fifo_csv_dumper_49,fifo_intf_49,cstatus_csv_dumper_49);
    fifo_csv_dumper_50 = new("./depth50.csv");
    cstatus_csv_dumper_50 = new("./chan_status50.csv");
    fifo_monitor_50 = new(fifo_csv_dumper_50,fifo_intf_50,cstatus_csv_dumper_50);
    fifo_csv_dumper_51 = new("./depth51.csv");
    cstatus_csv_dumper_51 = new("./chan_status51.csv");
    fifo_monitor_51 = new(fifo_csv_dumper_51,fifo_intf_51,cstatus_csv_dumper_51);
    fifo_csv_dumper_52 = new("./depth52.csv");
    cstatus_csv_dumper_52 = new("./chan_status52.csv");
    fifo_monitor_52 = new(fifo_csv_dumper_52,fifo_intf_52,cstatus_csv_dumper_52);
    fifo_csv_dumper_53 = new("./depth53.csv");
    cstatus_csv_dumper_53 = new("./chan_status53.csv");
    fifo_monitor_53 = new(fifo_csv_dumper_53,fifo_intf_53,cstatus_csv_dumper_53);
    fifo_csv_dumper_54 = new("./depth54.csv");
    cstatus_csv_dumper_54 = new("./chan_status54.csv");
    fifo_monitor_54 = new(fifo_csv_dumper_54,fifo_intf_54,cstatus_csv_dumper_54);
    fifo_csv_dumper_55 = new("./depth55.csv");
    cstatus_csv_dumper_55 = new("./chan_status55.csv");
    fifo_monitor_55 = new(fifo_csv_dumper_55,fifo_intf_55,cstatus_csv_dumper_55);
    fifo_csv_dumper_56 = new("./depth56.csv");
    cstatus_csv_dumper_56 = new("./chan_status56.csv");
    fifo_monitor_56 = new(fifo_csv_dumper_56,fifo_intf_56,cstatus_csv_dumper_56);
    fifo_csv_dumper_57 = new("./depth57.csv");
    cstatus_csv_dumper_57 = new("./chan_status57.csv");
    fifo_monitor_57 = new(fifo_csv_dumper_57,fifo_intf_57,cstatus_csv_dumper_57);
    fifo_csv_dumper_58 = new("./depth58.csv");
    cstatus_csv_dumper_58 = new("./chan_status58.csv");
    fifo_monitor_58 = new(fifo_csv_dumper_58,fifo_intf_58,cstatus_csv_dumper_58);
    fifo_csv_dumper_59 = new("./depth59.csv");
    cstatus_csv_dumper_59 = new("./chan_status59.csv");
    fifo_monitor_59 = new(fifo_csv_dumper_59,fifo_intf_59,cstatus_csv_dumper_59);
    fifo_csv_dumper_60 = new("./depth60.csv");
    cstatus_csv_dumper_60 = new("./chan_status60.csv");
    fifo_monitor_60 = new(fifo_csv_dumper_60,fifo_intf_60,cstatus_csv_dumper_60);
    fifo_csv_dumper_61 = new("./depth61.csv");
    cstatus_csv_dumper_61 = new("./chan_status61.csv");
    fifo_monitor_61 = new(fifo_csv_dumper_61,fifo_intf_61,cstatus_csv_dumper_61);
    fifo_csv_dumper_62 = new("./depth62.csv");
    cstatus_csv_dumper_62 = new("./chan_status62.csv");
    fifo_monitor_62 = new(fifo_csv_dumper_62,fifo_intf_62,cstatus_csv_dumper_62);
    fifo_csv_dumper_63 = new("./depth63.csv");
    cstatus_csv_dumper_63 = new("./chan_status63.csv");
    fifo_monitor_63 = new(fifo_csv_dumper_63,fifo_intf_63,cstatus_csv_dumper_63);
    fifo_csv_dumper_64 = new("./depth64.csv");
    cstatus_csv_dumper_64 = new("./chan_status64.csv");
    fifo_monitor_64 = new(fifo_csv_dumper_64,fifo_intf_64,cstatus_csv_dumper_64);
    fifo_csv_dumper_65 = new("./depth65.csv");
    cstatus_csv_dumper_65 = new("./chan_status65.csv");
    fifo_monitor_65 = new(fifo_csv_dumper_65,fifo_intf_65,cstatus_csv_dumper_65);
    fifo_csv_dumper_66 = new("./depth66.csv");
    cstatus_csv_dumper_66 = new("./chan_status66.csv");
    fifo_monitor_66 = new(fifo_csv_dumper_66,fifo_intf_66,cstatus_csv_dumper_66);
    fifo_csv_dumper_67 = new("./depth67.csv");
    cstatus_csv_dumper_67 = new("./chan_status67.csv");
    fifo_monitor_67 = new(fifo_csv_dumper_67,fifo_intf_67,cstatus_csv_dumper_67);
    fifo_csv_dumper_68 = new("./depth68.csv");
    cstatus_csv_dumper_68 = new("./chan_status68.csv");
    fifo_monitor_68 = new(fifo_csv_dumper_68,fifo_intf_68,cstatus_csv_dumper_68);
    fifo_csv_dumper_69 = new("./depth69.csv");
    cstatus_csv_dumper_69 = new("./chan_status69.csv");
    fifo_monitor_69 = new(fifo_csv_dumper_69,fifo_intf_69,cstatus_csv_dumper_69);
    fifo_csv_dumper_70 = new("./depth70.csv");
    cstatus_csv_dumper_70 = new("./chan_status70.csv");
    fifo_monitor_70 = new(fifo_csv_dumper_70,fifo_intf_70,cstatus_csv_dumper_70);
    fifo_csv_dumper_71 = new("./depth71.csv");
    cstatus_csv_dumper_71 = new("./chan_status71.csv");
    fifo_monitor_71 = new(fifo_csv_dumper_71,fifo_intf_71,cstatus_csv_dumper_71);
    fifo_csv_dumper_72 = new("./depth72.csv");
    cstatus_csv_dumper_72 = new("./chan_status72.csv");
    fifo_monitor_72 = new(fifo_csv_dumper_72,fifo_intf_72,cstatus_csv_dumper_72);
    fifo_csv_dumper_73 = new("./depth73.csv");
    cstatus_csv_dumper_73 = new("./chan_status73.csv");
    fifo_monitor_73 = new(fifo_csv_dumper_73,fifo_intf_73,cstatus_csv_dumper_73);
    fifo_csv_dumper_74 = new("./depth74.csv");
    cstatus_csv_dumper_74 = new("./chan_status74.csv");
    fifo_monitor_74 = new(fifo_csv_dumper_74,fifo_intf_74,cstatus_csv_dumper_74);
    fifo_csv_dumper_75 = new("./depth75.csv");
    cstatus_csv_dumper_75 = new("./chan_status75.csv");
    fifo_monitor_75 = new(fifo_csv_dumper_75,fifo_intf_75,cstatus_csv_dumper_75);
    fifo_csv_dumper_76 = new("./depth76.csv");
    cstatus_csv_dumper_76 = new("./chan_status76.csv");
    fifo_monitor_76 = new(fifo_csv_dumper_76,fifo_intf_76,cstatus_csv_dumper_76);
    fifo_csv_dumper_77 = new("./depth77.csv");
    cstatus_csv_dumper_77 = new("./chan_status77.csv");
    fifo_monitor_77 = new(fifo_csv_dumper_77,fifo_intf_77,cstatus_csv_dumper_77);
    fifo_csv_dumper_78 = new("./depth78.csv");
    cstatus_csv_dumper_78 = new("./chan_status78.csv");
    fifo_monitor_78 = new(fifo_csv_dumper_78,fifo_intf_78,cstatus_csv_dumper_78);
    fifo_csv_dumper_79 = new("./depth79.csv");
    cstatus_csv_dumper_79 = new("./chan_status79.csv");
    fifo_monitor_79 = new(fifo_csv_dumper_79,fifo_intf_79,cstatus_csv_dumper_79);
    fifo_csv_dumper_80 = new("./depth80.csv");
    cstatus_csv_dumper_80 = new("./chan_status80.csv");
    fifo_monitor_80 = new(fifo_csv_dumper_80,fifo_intf_80,cstatus_csv_dumper_80);
    fifo_csv_dumper_81 = new("./depth81.csv");
    cstatus_csv_dumper_81 = new("./chan_status81.csv");
    fifo_monitor_81 = new(fifo_csv_dumper_81,fifo_intf_81,cstatus_csv_dumper_81);
    fifo_csv_dumper_82 = new("./depth82.csv");
    cstatus_csv_dumper_82 = new("./chan_status82.csv");
    fifo_monitor_82 = new(fifo_csv_dumper_82,fifo_intf_82,cstatus_csv_dumper_82);
    fifo_csv_dumper_83 = new("./depth83.csv");
    cstatus_csv_dumper_83 = new("./chan_status83.csv");
    fifo_monitor_83 = new(fifo_csv_dumper_83,fifo_intf_83,cstatus_csv_dumper_83);
    fifo_csv_dumper_84 = new("./depth84.csv");
    cstatus_csv_dumper_84 = new("./chan_status84.csv");
    fifo_monitor_84 = new(fifo_csv_dumper_84,fifo_intf_84,cstatus_csv_dumper_84);
    fifo_csv_dumper_85 = new("./depth85.csv");
    cstatus_csv_dumper_85 = new("./chan_status85.csv");
    fifo_monitor_85 = new(fifo_csv_dumper_85,fifo_intf_85,cstatus_csv_dumper_85);
    fifo_csv_dumper_86 = new("./depth86.csv");
    cstatus_csv_dumper_86 = new("./chan_status86.csv");
    fifo_monitor_86 = new(fifo_csv_dumper_86,fifo_intf_86,cstatus_csv_dumper_86);
    fifo_csv_dumper_87 = new("./depth87.csv");
    cstatus_csv_dumper_87 = new("./chan_status87.csv");
    fifo_monitor_87 = new(fifo_csv_dumper_87,fifo_intf_87,cstatus_csv_dumper_87);
    fifo_csv_dumper_88 = new("./depth88.csv");
    cstatus_csv_dumper_88 = new("./chan_status88.csv");
    fifo_monitor_88 = new(fifo_csv_dumper_88,fifo_intf_88,cstatus_csv_dumper_88);
    fifo_csv_dumper_89 = new("./depth89.csv");
    cstatus_csv_dumper_89 = new("./chan_status89.csv");
    fifo_monitor_89 = new(fifo_csv_dumper_89,fifo_intf_89,cstatus_csv_dumper_89);
    fifo_csv_dumper_90 = new("./depth90.csv");
    cstatus_csv_dumper_90 = new("./chan_status90.csv");
    fifo_monitor_90 = new(fifo_csv_dumper_90,fifo_intf_90,cstatus_csv_dumper_90);
    fifo_csv_dumper_91 = new("./depth91.csv");
    cstatus_csv_dumper_91 = new("./chan_status91.csv");
    fifo_monitor_91 = new(fifo_csv_dumper_91,fifo_intf_91,cstatus_csv_dumper_91);
    fifo_csv_dumper_92 = new("./depth92.csv");
    cstatus_csv_dumper_92 = new("./chan_status92.csv");
    fifo_monitor_92 = new(fifo_csv_dumper_92,fifo_intf_92,cstatus_csv_dumper_92);
    fifo_csv_dumper_93 = new("./depth93.csv");
    cstatus_csv_dumper_93 = new("./chan_status93.csv");
    fifo_monitor_93 = new(fifo_csv_dumper_93,fifo_intf_93,cstatus_csv_dumper_93);
    fifo_csv_dumper_94 = new("./depth94.csv");
    cstatus_csv_dumper_94 = new("./chan_status94.csv");
    fifo_monitor_94 = new(fifo_csv_dumper_94,fifo_intf_94,cstatus_csv_dumper_94);
    fifo_csv_dumper_95 = new("./depth95.csv");
    cstatus_csv_dumper_95 = new("./chan_status95.csv");
    fifo_monitor_95 = new(fifo_csv_dumper_95,fifo_intf_95,cstatus_csv_dumper_95);
    fifo_csv_dumper_96 = new("./depth96.csv");
    cstatus_csv_dumper_96 = new("./chan_status96.csv");
    fifo_monitor_96 = new(fifo_csv_dumper_96,fifo_intf_96,cstatus_csv_dumper_96);
    fifo_csv_dumper_97 = new("./depth97.csv");
    cstatus_csv_dumper_97 = new("./chan_status97.csv");
    fifo_monitor_97 = new(fifo_csv_dumper_97,fifo_intf_97,cstatus_csv_dumper_97);
    fifo_csv_dumper_98 = new("./depth98.csv");
    cstatus_csv_dumper_98 = new("./chan_status98.csv");
    fifo_monitor_98 = new(fifo_csv_dumper_98,fifo_intf_98,cstatus_csv_dumper_98);
    fifo_csv_dumper_99 = new("./depth99.csv");
    cstatus_csv_dumper_99 = new("./chan_status99.csv");
    fifo_monitor_99 = new(fifo_csv_dumper_99,fifo_intf_99,cstatus_csv_dumper_99);
    fifo_csv_dumper_100 = new("./depth100.csv");
    cstatus_csv_dumper_100 = new("./chan_status100.csv");
    fifo_monitor_100 = new(fifo_csv_dumper_100,fifo_intf_100,cstatus_csv_dumper_100);
    fifo_csv_dumper_101 = new("./depth101.csv");
    cstatus_csv_dumper_101 = new("./chan_status101.csv");
    fifo_monitor_101 = new(fifo_csv_dumper_101,fifo_intf_101,cstatus_csv_dumper_101);
    fifo_csv_dumper_102 = new("./depth102.csv");
    cstatus_csv_dumper_102 = new("./chan_status102.csv");
    fifo_monitor_102 = new(fifo_csv_dumper_102,fifo_intf_102,cstatus_csv_dumper_102);
    fifo_csv_dumper_103 = new("./depth103.csv");
    cstatus_csv_dumper_103 = new("./chan_status103.csv");
    fifo_monitor_103 = new(fifo_csv_dumper_103,fifo_intf_103,cstatus_csv_dumper_103);
    fifo_csv_dumper_104 = new("./depth104.csv");
    cstatus_csv_dumper_104 = new("./chan_status104.csv");
    fifo_monitor_104 = new(fifo_csv_dumper_104,fifo_intf_104,cstatus_csv_dumper_104);
    fifo_csv_dumper_105 = new("./depth105.csv");
    cstatus_csv_dumper_105 = new("./chan_status105.csv");
    fifo_monitor_105 = new(fifo_csv_dumper_105,fifo_intf_105,cstatus_csv_dumper_105);
    fifo_csv_dumper_106 = new("./depth106.csv");
    cstatus_csv_dumper_106 = new("./chan_status106.csv");
    fifo_monitor_106 = new(fifo_csv_dumper_106,fifo_intf_106,cstatus_csv_dumper_106);
    fifo_csv_dumper_107 = new("./depth107.csv");
    cstatus_csv_dumper_107 = new("./chan_status107.csv");
    fifo_monitor_107 = new(fifo_csv_dumper_107,fifo_intf_107,cstatus_csv_dumper_107);
    fifo_csv_dumper_108 = new("./depth108.csv");
    cstatus_csv_dumper_108 = new("./chan_status108.csv");
    fifo_monitor_108 = new(fifo_csv_dumper_108,fifo_intf_108,cstatus_csv_dumper_108);
    fifo_csv_dumper_109 = new("./depth109.csv");
    cstatus_csv_dumper_109 = new("./chan_status109.csv");
    fifo_monitor_109 = new(fifo_csv_dumper_109,fifo_intf_109,cstatus_csv_dumper_109);
    fifo_csv_dumper_110 = new("./depth110.csv");
    cstatus_csv_dumper_110 = new("./chan_status110.csv");
    fifo_monitor_110 = new(fifo_csv_dumper_110,fifo_intf_110,cstatus_csv_dumper_110);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);




    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(fifo_monitor_18);
    sample_manager_inst.add_one_monitor(fifo_monitor_19);
    sample_manager_inst.add_one_monitor(fifo_monitor_20);
    sample_manager_inst.add_one_monitor(fifo_monitor_21);
    sample_manager_inst.add_one_monitor(fifo_monitor_22);
    sample_manager_inst.add_one_monitor(fifo_monitor_23);
    sample_manager_inst.add_one_monitor(fifo_monitor_24);
    sample_manager_inst.add_one_monitor(fifo_monitor_25);
    sample_manager_inst.add_one_monitor(fifo_monitor_26);
    sample_manager_inst.add_one_monitor(fifo_monitor_27);
    sample_manager_inst.add_one_monitor(fifo_monitor_28);
    sample_manager_inst.add_one_monitor(fifo_monitor_29);
    sample_manager_inst.add_one_monitor(fifo_monitor_30);
    sample_manager_inst.add_one_monitor(fifo_monitor_31);
    sample_manager_inst.add_one_monitor(fifo_monitor_32);
    sample_manager_inst.add_one_monitor(fifo_monitor_33);
    sample_manager_inst.add_one_monitor(fifo_monitor_34);
    sample_manager_inst.add_one_monitor(fifo_monitor_35);
    sample_manager_inst.add_one_monitor(fifo_monitor_36);
    sample_manager_inst.add_one_monitor(fifo_monitor_37);
    sample_manager_inst.add_one_monitor(fifo_monitor_38);
    sample_manager_inst.add_one_monitor(fifo_monitor_39);
    sample_manager_inst.add_one_monitor(fifo_monitor_40);
    sample_manager_inst.add_one_monitor(fifo_monitor_41);
    sample_manager_inst.add_one_monitor(fifo_monitor_42);
    sample_manager_inst.add_one_monitor(fifo_monitor_43);
    sample_manager_inst.add_one_monitor(fifo_monitor_44);
    sample_manager_inst.add_one_monitor(fifo_monitor_45);
    sample_manager_inst.add_one_monitor(fifo_monitor_46);
    sample_manager_inst.add_one_monitor(fifo_monitor_47);
    sample_manager_inst.add_one_monitor(fifo_monitor_48);
    sample_manager_inst.add_one_monitor(fifo_monitor_49);
    sample_manager_inst.add_one_monitor(fifo_monitor_50);
    sample_manager_inst.add_one_monitor(fifo_monitor_51);
    sample_manager_inst.add_one_monitor(fifo_monitor_52);
    sample_manager_inst.add_one_monitor(fifo_monitor_53);
    sample_manager_inst.add_one_monitor(fifo_monitor_54);
    sample_manager_inst.add_one_monitor(fifo_monitor_55);
    sample_manager_inst.add_one_monitor(fifo_monitor_56);
    sample_manager_inst.add_one_monitor(fifo_monitor_57);
    sample_manager_inst.add_one_monitor(fifo_monitor_58);
    sample_manager_inst.add_one_monitor(fifo_monitor_59);
    sample_manager_inst.add_one_monitor(fifo_monitor_60);
    sample_manager_inst.add_one_monitor(fifo_monitor_61);
    sample_manager_inst.add_one_monitor(fifo_monitor_62);
    sample_manager_inst.add_one_monitor(fifo_monitor_63);
    sample_manager_inst.add_one_monitor(fifo_monitor_64);
    sample_manager_inst.add_one_monitor(fifo_monitor_65);
    sample_manager_inst.add_one_monitor(fifo_monitor_66);
    sample_manager_inst.add_one_monitor(fifo_monitor_67);
    sample_manager_inst.add_one_monitor(fifo_monitor_68);
    sample_manager_inst.add_one_monitor(fifo_monitor_69);
    sample_manager_inst.add_one_monitor(fifo_monitor_70);
    sample_manager_inst.add_one_monitor(fifo_monitor_71);
    sample_manager_inst.add_one_monitor(fifo_monitor_72);
    sample_manager_inst.add_one_monitor(fifo_monitor_73);
    sample_manager_inst.add_one_monitor(fifo_monitor_74);
    sample_manager_inst.add_one_monitor(fifo_monitor_75);
    sample_manager_inst.add_one_monitor(fifo_monitor_76);
    sample_manager_inst.add_one_monitor(fifo_monitor_77);
    sample_manager_inst.add_one_monitor(fifo_monitor_78);
    sample_manager_inst.add_one_monitor(fifo_monitor_79);
    sample_manager_inst.add_one_monitor(fifo_monitor_80);
    sample_manager_inst.add_one_monitor(fifo_monitor_81);
    sample_manager_inst.add_one_monitor(fifo_monitor_82);
    sample_manager_inst.add_one_monitor(fifo_monitor_83);
    sample_manager_inst.add_one_monitor(fifo_monitor_84);
    sample_manager_inst.add_one_monitor(fifo_monitor_85);
    sample_manager_inst.add_one_monitor(fifo_monitor_86);
    sample_manager_inst.add_one_monitor(fifo_monitor_87);
    sample_manager_inst.add_one_monitor(fifo_monitor_88);
    sample_manager_inst.add_one_monitor(fifo_monitor_89);
    sample_manager_inst.add_one_monitor(fifo_monitor_90);
    sample_manager_inst.add_one_monitor(fifo_monitor_91);
    sample_manager_inst.add_one_monitor(fifo_monitor_92);
    sample_manager_inst.add_one_monitor(fifo_monitor_93);
    sample_manager_inst.add_one_monitor(fifo_monitor_94);
    sample_manager_inst.add_one_monitor(fifo_monitor_95);
    sample_manager_inst.add_one_monitor(fifo_monitor_96);
    sample_manager_inst.add_one_monitor(fifo_monitor_97);
    sample_manager_inst.add_one_monitor(fifo_monitor_98);
    sample_manager_inst.add_one_monitor(fifo_monitor_99);
    sample_manager_inst.add_one_monitor(fifo_monitor_100);
    sample_manager_inst.add_one_monitor(fifo_monitor_101);
    sample_manager_inst.add_one_monitor(fifo_monitor_102);
    sample_manager_inst.add_one_monitor(fifo_monitor_103);
    sample_manager_inst.add_one_monitor(fifo_monitor_104);
    sample_manager_inst.add_one_monitor(fifo_monitor_105);
    sample_manager_inst.add_one_monitor(fifo_monitor_106);
    sample_manager_inst.add_one_monitor(fifo_monitor_107);
    sample_manager_inst.add_one_monitor(fifo_monitor_108);
    sample_manager_inst.add_one_monitor(fifo_monitor_109);
    sample_manager_inst.add_one_monitor(fifo_monitor_110);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
